VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Integrated_bitcell_with_dummy_cells
  CLASS BLOCK ;
  FOREIGN Integrated_bitcell_with_dummy_cells ;
  ORIGIN 45.520 90.350 ;
  SIZE 191.920 BY 143.910 ;
  PIN PRE_SRAM
    ANTENNAGATEAREA 3.024000 ;
    PORT
      LAYER met1 ;
        RECT 4.340 50.140 4.670 50.190 ;
        RECT 5.210 50.140 5.540 50.190 ;
        RECT 6.080 50.140 6.410 50.190 ;
        RECT 10.090 50.140 10.420 50.190 ;
        RECT 10.960 50.140 11.290 50.190 ;
        RECT 11.830 50.140 12.160 50.190 ;
        RECT 15.840 50.140 16.170 50.190 ;
        RECT 16.710 50.140 17.040 50.190 ;
        RECT 17.580 50.140 17.910 50.190 ;
        RECT 21.590 50.140 21.920 50.190 ;
        RECT 22.460 50.140 22.790 50.190 ;
        RECT 23.330 50.140 23.660 50.190 ;
        RECT 27.340 50.140 27.670 50.190 ;
        RECT 28.210 50.140 28.540 50.190 ;
        RECT 29.080 50.140 29.410 50.190 ;
        RECT 33.090 50.140 33.420 50.190 ;
        RECT 33.960 50.140 34.290 50.190 ;
        RECT 34.830 50.140 35.160 50.190 ;
        RECT 38.840 50.140 39.170 50.190 ;
        RECT 39.710 50.140 40.040 50.190 ;
        RECT 40.580 50.140 40.910 50.190 ;
        RECT 44.590 50.140 44.920 50.190 ;
        RECT 45.460 50.140 45.790 50.190 ;
        RECT 46.330 50.140 46.660 50.190 ;
        RECT 50.340 50.140 50.670 50.190 ;
        RECT 51.210 50.140 51.540 50.190 ;
        RECT 52.080 50.140 52.410 50.190 ;
        RECT 56.090 50.140 56.420 50.190 ;
        RECT 56.960 50.140 57.290 50.190 ;
        RECT 57.830 50.140 58.160 50.190 ;
        RECT 61.840 50.140 62.170 50.190 ;
        RECT 62.710 50.140 63.040 50.190 ;
        RECT 63.580 50.140 63.910 50.190 ;
        RECT 67.590 50.140 67.920 50.190 ;
        RECT 68.460 50.140 68.790 50.190 ;
        RECT 69.330 50.140 69.660 50.190 ;
        RECT 73.340 50.140 73.670 50.190 ;
        RECT 74.210 50.140 74.540 50.190 ;
        RECT 75.080 50.140 75.410 50.190 ;
        RECT 79.090 50.140 79.420 50.190 ;
        RECT 79.960 50.140 80.290 50.190 ;
        RECT 80.830 50.140 81.160 50.190 ;
        RECT 84.840 50.140 85.170 50.190 ;
        RECT 85.710 50.140 86.040 50.190 ;
        RECT 86.580 50.140 86.910 50.190 ;
        RECT 90.590 50.140 90.920 50.190 ;
        RECT 91.460 50.140 91.790 50.190 ;
        RECT 92.330 50.140 92.660 50.190 ;
        RECT -45.490 50.000 94.660 50.140 ;
        RECT 4.340 49.960 4.670 50.000 ;
        RECT 5.210 49.960 5.540 50.000 ;
        RECT 6.080 49.960 6.410 50.000 ;
        RECT 10.090 49.960 10.420 50.000 ;
        RECT 10.960 49.960 11.290 50.000 ;
        RECT 11.830 49.960 12.160 50.000 ;
        RECT 15.840 49.960 16.170 50.000 ;
        RECT 16.710 49.960 17.040 50.000 ;
        RECT 17.580 49.960 17.910 50.000 ;
        RECT 21.590 49.960 21.920 50.000 ;
        RECT 22.460 49.960 22.790 50.000 ;
        RECT 23.330 49.960 23.660 50.000 ;
        RECT 27.340 49.960 27.670 50.000 ;
        RECT 28.210 49.960 28.540 50.000 ;
        RECT 29.080 49.960 29.410 50.000 ;
        RECT 33.090 49.960 33.420 50.000 ;
        RECT 33.960 49.960 34.290 50.000 ;
        RECT 34.830 49.960 35.160 50.000 ;
        RECT 38.840 49.960 39.170 50.000 ;
        RECT 39.710 49.960 40.040 50.000 ;
        RECT 40.580 49.960 40.910 50.000 ;
        RECT 44.590 49.960 44.920 50.000 ;
        RECT 45.460 49.960 45.790 50.000 ;
        RECT 46.330 49.960 46.660 50.000 ;
        RECT 50.340 49.960 50.670 50.000 ;
        RECT 51.210 49.960 51.540 50.000 ;
        RECT 52.080 49.960 52.410 50.000 ;
        RECT 56.090 49.960 56.420 50.000 ;
        RECT 56.960 49.960 57.290 50.000 ;
        RECT 57.830 49.960 58.160 50.000 ;
        RECT 61.840 49.960 62.170 50.000 ;
        RECT 62.710 49.960 63.040 50.000 ;
        RECT 63.580 49.960 63.910 50.000 ;
        RECT 67.590 49.960 67.920 50.000 ;
        RECT 68.460 49.960 68.790 50.000 ;
        RECT 69.330 49.960 69.660 50.000 ;
        RECT 73.340 49.960 73.670 50.000 ;
        RECT 74.210 49.960 74.540 50.000 ;
        RECT 75.080 49.960 75.410 50.000 ;
        RECT 79.090 49.960 79.420 50.000 ;
        RECT 79.960 49.960 80.290 50.000 ;
        RECT 80.830 49.960 81.160 50.000 ;
        RECT 84.840 49.960 85.170 50.000 ;
        RECT 85.710 49.960 86.040 50.000 ;
        RECT 86.580 49.960 86.910 50.000 ;
        RECT 90.590 49.960 90.920 50.000 ;
        RECT 91.460 49.960 91.790 50.000 ;
        RECT 92.330 49.960 92.660 50.000 ;
    END
  END PRE_SRAM
  PIN RWL[0]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 37.550 2.760 37.620 ;
        RECT 8.210 37.550 8.510 37.620 ;
        RECT 13.960 37.550 14.260 37.620 ;
        RECT 19.710 37.550 20.010 37.620 ;
        RECT 25.460 37.550 25.760 37.620 ;
        RECT 31.210 37.550 31.510 37.620 ;
        RECT 36.960 37.550 37.260 37.620 ;
        RECT 42.710 37.550 43.010 37.620 ;
        RECT 48.460 37.550 48.760 37.620 ;
        RECT 54.210 37.550 54.510 37.620 ;
        RECT 59.960 37.550 60.260 37.620 ;
        RECT 65.710 37.550 66.010 37.620 ;
        RECT 71.460 37.550 71.760 37.620 ;
        RECT 77.210 37.550 77.510 37.620 ;
        RECT 82.960 37.550 83.260 37.620 ;
        RECT 88.710 37.550 89.010 37.620 ;
        RECT -45.490 37.410 94.660 37.550 ;
        RECT 2.460 37.330 2.760 37.410 ;
        RECT 8.210 37.330 8.510 37.410 ;
        RECT 13.960 37.330 14.260 37.410 ;
        RECT 19.710 37.330 20.010 37.410 ;
        RECT 25.460 37.330 25.760 37.410 ;
        RECT 31.210 37.330 31.510 37.410 ;
        RECT 36.960 37.330 37.260 37.410 ;
        RECT 42.710 37.330 43.010 37.410 ;
        RECT 48.460 37.330 48.760 37.410 ;
        RECT 54.210 37.330 54.510 37.410 ;
        RECT 59.960 37.330 60.260 37.410 ;
        RECT 65.710 37.330 66.010 37.410 ;
        RECT 71.460 37.330 71.760 37.410 ;
        RECT 77.210 37.330 77.510 37.410 ;
        RECT 82.960 37.330 83.260 37.410 ;
        RECT 88.710 37.330 89.010 37.410 ;
    END
  END RWL[0]
  PIN WWL[0]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 37.150 4.730 37.270 ;
        RECT 10.190 37.150 10.480 37.270 ;
        RECT 15.940 37.150 16.230 37.270 ;
        RECT 21.690 37.150 21.980 37.270 ;
        RECT 27.440 37.150 27.730 37.270 ;
        RECT 33.190 37.150 33.480 37.270 ;
        RECT 38.940 37.150 39.230 37.270 ;
        RECT 44.690 37.150 44.980 37.270 ;
        RECT 50.440 37.150 50.730 37.270 ;
        RECT 56.190 37.150 56.480 37.270 ;
        RECT 61.940 37.150 62.230 37.270 ;
        RECT 67.690 37.150 67.980 37.270 ;
        RECT 73.440 37.150 73.730 37.270 ;
        RECT 79.190 37.150 79.480 37.270 ;
        RECT 84.940 37.150 85.230 37.270 ;
        RECT 90.690 37.150 90.980 37.270 ;
        RECT -45.490 37.010 94.660 37.150 ;
        RECT 6.050 36.890 6.340 37.010 ;
        RECT 11.800 36.890 12.090 37.010 ;
        RECT 17.550 36.890 17.840 37.010 ;
        RECT 23.300 36.890 23.590 37.010 ;
        RECT 29.050 36.890 29.340 37.010 ;
        RECT 34.800 36.890 35.090 37.010 ;
        RECT 40.550 36.890 40.840 37.010 ;
        RECT 46.300 36.890 46.590 37.010 ;
        RECT 52.050 36.890 52.340 37.010 ;
        RECT 57.800 36.890 58.090 37.010 ;
        RECT 63.550 36.890 63.840 37.010 ;
        RECT 69.300 36.890 69.590 37.010 ;
        RECT 75.050 36.890 75.340 37.010 ;
        RECT 80.800 36.890 81.090 37.010 ;
        RECT 86.550 36.890 86.840 37.010 ;
        RECT 92.300 36.890 92.590 37.010 ;
    END
  END WWL[0]
  PIN RWLB[0]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 36.740 8.310 36.840 ;
        RECT 13.760 36.740 14.060 36.840 ;
        RECT 19.510 36.740 19.810 36.840 ;
        RECT 25.260 36.740 25.560 36.840 ;
        RECT 31.010 36.740 31.310 36.840 ;
        RECT 36.760 36.740 37.060 36.840 ;
        RECT 42.510 36.740 42.810 36.840 ;
        RECT 48.260 36.740 48.560 36.840 ;
        RECT 54.010 36.740 54.310 36.840 ;
        RECT 59.760 36.740 60.060 36.840 ;
        RECT 65.510 36.740 65.810 36.840 ;
        RECT 71.260 36.740 71.560 36.840 ;
        RECT 77.010 36.740 77.310 36.840 ;
        RECT 82.760 36.740 83.060 36.840 ;
        RECT 88.510 36.740 88.810 36.840 ;
        RECT 94.260 36.740 94.560 36.840 ;
        RECT -45.490 36.600 94.660 36.740 ;
        RECT 8.010 36.510 8.310 36.600 ;
        RECT 13.760 36.510 14.060 36.600 ;
        RECT 19.510 36.510 19.810 36.600 ;
        RECT 25.260 36.510 25.560 36.600 ;
        RECT 31.010 36.510 31.310 36.600 ;
        RECT 36.760 36.510 37.060 36.600 ;
        RECT 42.510 36.510 42.810 36.600 ;
        RECT 48.260 36.510 48.560 36.600 ;
        RECT 54.010 36.510 54.310 36.600 ;
        RECT 59.760 36.510 60.060 36.600 ;
        RECT 65.510 36.510 65.810 36.600 ;
        RECT 71.260 36.510 71.560 36.600 ;
        RECT 77.010 36.510 77.310 36.600 ;
        RECT 82.760 36.510 83.060 36.600 ;
        RECT 88.510 36.510 88.810 36.600 ;
        RECT 94.260 36.510 94.560 36.600 ;
    END
  END RWLB[0]
  PIN RWL[1]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 35.140 2.760 35.210 ;
        RECT 8.210 35.140 8.510 35.210 ;
        RECT 13.960 35.140 14.260 35.210 ;
        RECT 19.710 35.140 20.010 35.210 ;
        RECT 25.460 35.140 25.760 35.210 ;
        RECT 31.210 35.140 31.510 35.210 ;
        RECT 36.960 35.140 37.260 35.210 ;
        RECT 42.710 35.140 43.010 35.210 ;
        RECT 48.460 35.140 48.760 35.210 ;
        RECT 54.210 35.140 54.510 35.210 ;
        RECT 59.960 35.140 60.260 35.210 ;
        RECT 65.710 35.140 66.010 35.210 ;
        RECT 71.460 35.140 71.760 35.210 ;
        RECT 77.210 35.140 77.510 35.210 ;
        RECT 82.960 35.140 83.260 35.210 ;
        RECT 88.710 35.140 89.010 35.210 ;
        RECT -45.490 35.000 94.660 35.140 ;
        RECT 2.460 34.920 2.760 35.000 ;
        RECT 8.210 34.920 8.510 35.000 ;
        RECT 13.960 34.920 14.260 35.000 ;
        RECT 19.710 34.920 20.010 35.000 ;
        RECT 25.460 34.920 25.760 35.000 ;
        RECT 31.210 34.920 31.510 35.000 ;
        RECT 36.960 34.920 37.260 35.000 ;
        RECT 42.710 34.920 43.010 35.000 ;
        RECT 48.460 34.920 48.760 35.000 ;
        RECT 54.210 34.920 54.510 35.000 ;
        RECT 59.960 34.920 60.260 35.000 ;
        RECT 65.710 34.920 66.010 35.000 ;
        RECT 71.460 34.920 71.760 35.000 ;
        RECT 77.210 34.920 77.510 35.000 ;
        RECT 82.960 34.920 83.260 35.000 ;
        RECT 88.710 34.920 89.010 35.000 ;
    END
  END RWL[1]
  PIN WWL[1]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 34.740 4.730 34.860 ;
        RECT 10.190 34.740 10.480 34.860 ;
        RECT 15.940 34.740 16.230 34.860 ;
        RECT 21.690 34.740 21.980 34.860 ;
        RECT 27.440 34.740 27.730 34.860 ;
        RECT 33.190 34.740 33.480 34.860 ;
        RECT 38.940 34.740 39.230 34.860 ;
        RECT 44.690 34.740 44.980 34.860 ;
        RECT 50.440 34.740 50.730 34.860 ;
        RECT 56.190 34.740 56.480 34.860 ;
        RECT 61.940 34.740 62.230 34.860 ;
        RECT 67.690 34.740 67.980 34.860 ;
        RECT 73.440 34.740 73.730 34.860 ;
        RECT 79.190 34.740 79.480 34.860 ;
        RECT 84.940 34.740 85.230 34.860 ;
        RECT 90.690 34.740 90.980 34.860 ;
        RECT -45.490 34.600 94.660 34.740 ;
        RECT 6.050 34.480 6.340 34.600 ;
        RECT 11.800 34.480 12.090 34.600 ;
        RECT 17.550 34.480 17.840 34.600 ;
        RECT 23.300 34.480 23.590 34.600 ;
        RECT 29.050 34.480 29.340 34.600 ;
        RECT 34.800 34.480 35.090 34.600 ;
        RECT 40.550 34.480 40.840 34.600 ;
        RECT 46.300 34.480 46.590 34.600 ;
        RECT 52.050 34.480 52.340 34.600 ;
        RECT 57.800 34.480 58.090 34.600 ;
        RECT 63.550 34.480 63.840 34.600 ;
        RECT 69.300 34.480 69.590 34.600 ;
        RECT 75.050 34.480 75.340 34.600 ;
        RECT 80.800 34.480 81.090 34.600 ;
        RECT 86.550 34.480 86.840 34.600 ;
        RECT 92.300 34.480 92.590 34.600 ;
    END
  END WWL[1]
  PIN RWLB[1]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 34.330 8.310 34.430 ;
        RECT 13.760 34.330 14.060 34.430 ;
        RECT 19.510 34.330 19.810 34.430 ;
        RECT 25.260 34.330 25.560 34.430 ;
        RECT 31.010 34.330 31.310 34.430 ;
        RECT 36.760 34.330 37.060 34.430 ;
        RECT 42.510 34.330 42.810 34.430 ;
        RECT 48.260 34.330 48.560 34.430 ;
        RECT 54.010 34.330 54.310 34.430 ;
        RECT 59.760 34.330 60.060 34.430 ;
        RECT 65.510 34.330 65.810 34.430 ;
        RECT 71.260 34.330 71.560 34.430 ;
        RECT 77.010 34.330 77.310 34.430 ;
        RECT 82.760 34.330 83.060 34.430 ;
        RECT 88.510 34.330 88.810 34.430 ;
        RECT 94.260 34.330 94.560 34.430 ;
        RECT -45.490 34.190 94.660 34.330 ;
        RECT 8.010 34.100 8.310 34.190 ;
        RECT 13.760 34.100 14.060 34.190 ;
        RECT 19.510 34.100 19.810 34.190 ;
        RECT 25.260 34.100 25.560 34.190 ;
        RECT 31.010 34.100 31.310 34.190 ;
        RECT 36.760 34.100 37.060 34.190 ;
        RECT 42.510 34.100 42.810 34.190 ;
        RECT 48.260 34.100 48.560 34.190 ;
        RECT 54.010 34.100 54.310 34.190 ;
        RECT 59.760 34.100 60.060 34.190 ;
        RECT 65.510 34.100 65.810 34.190 ;
        RECT 71.260 34.100 71.560 34.190 ;
        RECT 77.010 34.100 77.310 34.190 ;
        RECT 82.760 34.100 83.060 34.190 ;
        RECT 88.510 34.100 88.810 34.190 ;
        RECT 94.260 34.100 94.560 34.190 ;
    END
  END RWLB[1]
  PIN RWL[2]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 32.730 2.760 32.800 ;
        RECT 8.210 32.730 8.510 32.800 ;
        RECT 13.960 32.730 14.260 32.800 ;
        RECT 19.710 32.730 20.010 32.800 ;
        RECT 25.460 32.730 25.760 32.800 ;
        RECT 31.210 32.730 31.510 32.800 ;
        RECT 36.960 32.730 37.260 32.800 ;
        RECT 42.710 32.730 43.010 32.800 ;
        RECT 48.460 32.730 48.760 32.800 ;
        RECT 54.210 32.730 54.510 32.800 ;
        RECT 59.960 32.730 60.260 32.800 ;
        RECT 65.710 32.730 66.010 32.800 ;
        RECT 71.460 32.730 71.760 32.800 ;
        RECT 77.210 32.730 77.510 32.800 ;
        RECT 82.960 32.730 83.260 32.800 ;
        RECT 88.710 32.730 89.010 32.800 ;
        RECT -45.490 32.590 94.660 32.730 ;
        RECT 2.460 32.510 2.760 32.590 ;
        RECT 8.210 32.510 8.510 32.590 ;
        RECT 13.960 32.510 14.260 32.590 ;
        RECT 19.710 32.510 20.010 32.590 ;
        RECT 25.460 32.510 25.760 32.590 ;
        RECT 31.210 32.510 31.510 32.590 ;
        RECT 36.960 32.510 37.260 32.590 ;
        RECT 42.710 32.510 43.010 32.590 ;
        RECT 48.460 32.510 48.760 32.590 ;
        RECT 54.210 32.510 54.510 32.590 ;
        RECT 59.960 32.510 60.260 32.590 ;
        RECT 65.710 32.510 66.010 32.590 ;
        RECT 71.460 32.510 71.760 32.590 ;
        RECT 77.210 32.510 77.510 32.590 ;
        RECT 82.960 32.510 83.260 32.590 ;
        RECT 88.710 32.510 89.010 32.590 ;
    END
  END RWL[2]
  PIN WWL[2]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 32.330 4.730 32.450 ;
        RECT 10.190 32.330 10.480 32.450 ;
        RECT 15.940 32.330 16.230 32.450 ;
        RECT 21.690 32.330 21.980 32.450 ;
        RECT 27.440 32.330 27.730 32.450 ;
        RECT 33.190 32.330 33.480 32.450 ;
        RECT 38.940 32.330 39.230 32.450 ;
        RECT 44.690 32.330 44.980 32.450 ;
        RECT 50.440 32.330 50.730 32.450 ;
        RECT 56.190 32.330 56.480 32.450 ;
        RECT 61.940 32.330 62.230 32.450 ;
        RECT 67.690 32.330 67.980 32.450 ;
        RECT 73.440 32.330 73.730 32.450 ;
        RECT 79.190 32.330 79.480 32.450 ;
        RECT 84.940 32.330 85.230 32.450 ;
        RECT 90.690 32.330 90.980 32.450 ;
        RECT -45.490 32.190 94.660 32.330 ;
        RECT 6.050 32.070 6.340 32.190 ;
        RECT 11.800 32.070 12.090 32.190 ;
        RECT 17.550 32.070 17.840 32.190 ;
        RECT 23.300 32.070 23.590 32.190 ;
        RECT 29.050 32.070 29.340 32.190 ;
        RECT 34.800 32.070 35.090 32.190 ;
        RECT 40.550 32.070 40.840 32.190 ;
        RECT 46.300 32.070 46.590 32.190 ;
        RECT 52.050 32.070 52.340 32.190 ;
        RECT 57.800 32.070 58.090 32.190 ;
        RECT 63.550 32.070 63.840 32.190 ;
        RECT 69.300 32.070 69.590 32.190 ;
        RECT 75.050 32.070 75.340 32.190 ;
        RECT 80.800 32.070 81.090 32.190 ;
        RECT 86.550 32.070 86.840 32.190 ;
        RECT 92.300 32.070 92.590 32.190 ;
    END
  END WWL[2]
  PIN RWLB[2]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 31.920 8.310 32.020 ;
        RECT 13.760 31.920 14.060 32.020 ;
        RECT 19.510 31.920 19.810 32.020 ;
        RECT 25.260 31.920 25.560 32.020 ;
        RECT 31.010 31.920 31.310 32.020 ;
        RECT 36.760 31.920 37.060 32.020 ;
        RECT 42.510 31.920 42.810 32.020 ;
        RECT 48.260 31.920 48.560 32.020 ;
        RECT 54.010 31.920 54.310 32.020 ;
        RECT 59.760 31.920 60.060 32.020 ;
        RECT 65.510 31.920 65.810 32.020 ;
        RECT 71.260 31.920 71.560 32.020 ;
        RECT 77.010 31.920 77.310 32.020 ;
        RECT 82.760 31.920 83.060 32.020 ;
        RECT 88.510 31.920 88.810 32.020 ;
        RECT 94.260 31.920 94.560 32.020 ;
        RECT -45.490 31.780 94.660 31.920 ;
        RECT 8.010 31.690 8.310 31.780 ;
        RECT 13.760 31.690 14.060 31.780 ;
        RECT 19.510 31.690 19.810 31.780 ;
        RECT 25.260 31.690 25.560 31.780 ;
        RECT 31.010 31.690 31.310 31.780 ;
        RECT 36.760 31.690 37.060 31.780 ;
        RECT 42.510 31.690 42.810 31.780 ;
        RECT 48.260 31.690 48.560 31.780 ;
        RECT 54.010 31.690 54.310 31.780 ;
        RECT 59.760 31.690 60.060 31.780 ;
        RECT 65.510 31.690 65.810 31.780 ;
        RECT 71.260 31.690 71.560 31.780 ;
        RECT 77.010 31.690 77.310 31.780 ;
        RECT 82.760 31.690 83.060 31.780 ;
        RECT 88.510 31.690 88.810 31.780 ;
        RECT 94.260 31.690 94.560 31.780 ;
    END
  END RWLB[2]
  PIN RWL[3]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 30.320 2.760 30.390 ;
        RECT 8.210 30.320 8.510 30.390 ;
        RECT 13.960 30.320 14.260 30.390 ;
        RECT 19.710 30.320 20.010 30.390 ;
        RECT 25.460 30.320 25.760 30.390 ;
        RECT 31.210 30.320 31.510 30.390 ;
        RECT 36.960 30.320 37.260 30.390 ;
        RECT 42.710 30.320 43.010 30.390 ;
        RECT 48.460 30.320 48.760 30.390 ;
        RECT 54.210 30.320 54.510 30.390 ;
        RECT 59.960 30.320 60.260 30.390 ;
        RECT 65.710 30.320 66.010 30.390 ;
        RECT 71.460 30.320 71.760 30.390 ;
        RECT 77.210 30.320 77.510 30.390 ;
        RECT 82.960 30.320 83.260 30.390 ;
        RECT 88.710 30.320 89.010 30.390 ;
        RECT -45.490 30.180 94.660 30.320 ;
        RECT 2.460 30.100 2.760 30.180 ;
        RECT 8.210 30.100 8.510 30.180 ;
        RECT 13.960 30.100 14.260 30.180 ;
        RECT 19.710 30.100 20.010 30.180 ;
        RECT 25.460 30.100 25.760 30.180 ;
        RECT 31.210 30.100 31.510 30.180 ;
        RECT 36.960 30.100 37.260 30.180 ;
        RECT 42.710 30.100 43.010 30.180 ;
        RECT 48.460 30.100 48.760 30.180 ;
        RECT 54.210 30.100 54.510 30.180 ;
        RECT 59.960 30.100 60.260 30.180 ;
        RECT 65.710 30.100 66.010 30.180 ;
        RECT 71.460 30.100 71.760 30.180 ;
        RECT 77.210 30.100 77.510 30.180 ;
        RECT 82.960 30.100 83.260 30.180 ;
        RECT 88.710 30.100 89.010 30.180 ;
    END
  END RWL[3]
  PIN WWL[3]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 29.920 4.730 30.040 ;
        RECT 10.190 29.920 10.480 30.040 ;
        RECT 15.940 29.920 16.230 30.040 ;
        RECT 21.690 29.920 21.980 30.040 ;
        RECT 27.440 29.920 27.730 30.040 ;
        RECT 33.190 29.920 33.480 30.040 ;
        RECT 38.940 29.920 39.230 30.040 ;
        RECT 44.690 29.920 44.980 30.040 ;
        RECT 50.440 29.920 50.730 30.040 ;
        RECT 56.190 29.920 56.480 30.040 ;
        RECT 61.940 29.920 62.230 30.040 ;
        RECT 67.690 29.920 67.980 30.040 ;
        RECT 73.440 29.920 73.730 30.040 ;
        RECT 79.190 29.920 79.480 30.040 ;
        RECT 84.940 29.920 85.230 30.040 ;
        RECT 90.690 29.920 90.980 30.040 ;
        RECT -45.490 29.780 94.660 29.920 ;
        RECT 6.050 29.660 6.340 29.780 ;
        RECT 11.800 29.660 12.090 29.780 ;
        RECT 17.550 29.660 17.840 29.780 ;
        RECT 23.300 29.660 23.590 29.780 ;
        RECT 29.050 29.660 29.340 29.780 ;
        RECT 34.800 29.660 35.090 29.780 ;
        RECT 40.550 29.660 40.840 29.780 ;
        RECT 46.300 29.660 46.590 29.780 ;
        RECT 52.050 29.660 52.340 29.780 ;
        RECT 57.800 29.660 58.090 29.780 ;
        RECT 63.550 29.660 63.840 29.780 ;
        RECT 69.300 29.660 69.590 29.780 ;
        RECT 75.050 29.660 75.340 29.780 ;
        RECT 80.800 29.660 81.090 29.780 ;
        RECT 86.550 29.660 86.840 29.780 ;
        RECT 92.300 29.660 92.590 29.780 ;
    END
  END WWL[3]
  PIN RWLB[3]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 29.510 8.310 29.610 ;
        RECT 13.760 29.510 14.060 29.610 ;
        RECT 19.510 29.510 19.810 29.610 ;
        RECT 25.260 29.510 25.560 29.610 ;
        RECT 31.010 29.510 31.310 29.610 ;
        RECT 36.760 29.510 37.060 29.610 ;
        RECT 42.510 29.510 42.810 29.610 ;
        RECT 48.260 29.510 48.560 29.610 ;
        RECT 54.010 29.510 54.310 29.610 ;
        RECT 59.760 29.510 60.060 29.610 ;
        RECT 65.510 29.510 65.810 29.610 ;
        RECT 71.260 29.510 71.560 29.610 ;
        RECT 77.010 29.510 77.310 29.610 ;
        RECT 82.760 29.510 83.060 29.610 ;
        RECT 88.510 29.510 88.810 29.610 ;
        RECT 94.260 29.510 94.560 29.610 ;
        RECT -45.490 29.370 94.660 29.510 ;
        RECT 8.010 29.280 8.310 29.370 ;
        RECT 13.760 29.280 14.060 29.370 ;
        RECT 19.510 29.280 19.810 29.370 ;
        RECT 25.260 29.280 25.560 29.370 ;
        RECT 31.010 29.280 31.310 29.370 ;
        RECT 36.760 29.280 37.060 29.370 ;
        RECT 42.510 29.280 42.810 29.370 ;
        RECT 48.260 29.280 48.560 29.370 ;
        RECT 54.010 29.280 54.310 29.370 ;
        RECT 59.760 29.280 60.060 29.370 ;
        RECT 65.510 29.280 65.810 29.370 ;
        RECT 71.260 29.280 71.560 29.370 ;
        RECT 77.010 29.280 77.310 29.370 ;
        RECT 82.760 29.280 83.060 29.370 ;
        RECT 88.510 29.280 88.810 29.370 ;
        RECT 94.260 29.280 94.560 29.370 ;
    END
  END RWLB[3]
  PIN RWL[4]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 27.510 2.760 27.570 ;
        RECT 8.210 27.510 8.510 27.570 ;
        RECT 13.960 27.510 14.260 27.570 ;
        RECT 19.710 27.510 20.010 27.570 ;
        RECT 25.460 27.510 25.760 27.570 ;
        RECT 31.210 27.510 31.510 27.570 ;
        RECT 36.960 27.510 37.260 27.570 ;
        RECT 42.710 27.510 43.010 27.570 ;
        RECT 48.460 27.510 48.760 27.570 ;
        RECT 54.210 27.510 54.510 27.570 ;
        RECT 59.960 27.510 60.260 27.570 ;
        RECT 65.710 27.510 66.010 27.570 ;
        RECT 71.460 27.510 71.760 27.570 ;
        RECT 77.210 27.510 77.510 27.570 ;
        RECT 82.960 27.510 83.260 27.570 ;
        RECT 88.710 27.510 89.010 27.570 ;
        RECT -45.490 27.370 94.660 27.510 ;
        RECT 2.460 27.290 2.760 27.370 ;
        RECT 8.210 27.290 8.510 27.370 ;
        RECT 13.960 27.290 14.260 27.370 ;
        RECT 19.710 27.290 20.010 27.370 ;
        RECT 25.460 27.290 25.760 27.370 ;
        RECT 31.210 27.290 31.510 27.370 ;
        RECT 36.960 27.290 37.260 27.370 ;
        RECT 42.710 27.290 43.010 27.370 ;
        RECT 48.460 27.290 48.760 27.370 ;
        RECT 54.210 27.290 54.510 27.370 ;
        RECT 59.960 27.290 60.260 27.370 ;
        RECT 65.710 27.290 66.010 27.370 ;
        RECT 71.460 27.290 71.760 27.370 ;
        RECT 77.210 27.290 77.510 27.370 ;
        RECT 82.960 27.290 83.260 27.370 ;
        RECT 88.710 27.290 89.010 27.370 ;
    END
  END RWL[4]
  PIN WWL[4]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 27.110 4.730 27.230 ;
        RECT 10.190 27.110 10.480 27.230 ;
        RECT 15.940 27.110 16.230 27.230 ;
        RECT 21.690 27.110 21.980 27.230 ;
        RECT 27.440 27.110 27.730 27.230 ;
        RECT 33.190 27.110 33.480 27.230 ;
        RECT 38.940 27.110 39.230 27.230 ;
        RECT 44.690 27.110 44.980 27.230 ;
        RECT 50.440 27.110 50.730 27.230 ;
        RECT 56.190 27.110 56.480 27.230 ;
        RECT 61.940 27.110 62.230 27.230 ;
        RECT 67.690 27.110 67.980 27.230 ;
        RECT 73.440 27.110 73.730 27.230 ;
        RECT 79.190 27.110 79.480 27.230 ;
        RECT 84.940 27.110 85.230 27.230 ;
        RECT 90.690 27.110 90.980 27.230 ;
        RECT -45.490 26.970 94.660 27.110 ;
        RECT 6.050 26.850 6.340 26.970 ;
        RECT 11.800 26.850 12.090 26.970 ;
        RECT 17.550 26.850 17.840 26.970 ;
        RECT 23.300 26.850 23.590 26.970 ;
        RECT 29.050 26.850 29.340 26.970 ;
        RECT 34.800 26.850 35.090 26.970 ;
        RECT 40.550 26.850 40.840 26.970 ;
        RECT 46.300 26.850 46.590 26.970 ;
        RECT 52.050 26.850 52.340 26.970 ;
        RECT 57.800 26.850 58.090 26.970 ;
        RECT 63.550 26.850 63.840 26.970 ;
        RECT 69.300 26.850 69.590 26.970 ;
        RECT 75.050 26.850 75.340 26.970 ;
        RECT 80.800 26.850 81.090 26.970 ;
        RECT 86.550 26.850 86.840 26.970 ;
        RECT 92.300 26.850 92.590 26.970 ;
    END
  END WWL[4]
  PIN RWLB[4]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 26.700 8.310 26.800 ;
        RECT 13.760 26.700 14.060 26.800 ;
        RECT 19.510 26.700 19.810 26.800 ;
        RECT 25.260 26.700 25.560 26.800 ;
        RECT 31.010 26.700 31.310 26.800 ;
        RECT 36.760 26.700 37.060 26.800 ;
        RECT 42.510 26.700 42.810 26.800 ;
        RECT 48.260 26.700 48.560 26.800 ;
        RECT 54.010 26.700 54.310 26.800 ;
        RECT 59.760 26.700 60.060 26.800 ;
        RECT 65.510 26.700 65.810 26.800 ;
        RECT 71.260 26.700 71.560 26.800 ;
        RECT 77.010 26.700 77.310 26.800 ;
        RECT 82.760 26.700 83.060 26.800 ;
        RECT 88.510 26.700 88.810 26.800 ;
        RECT 94.260 26.700 94.560 26.800 ;
        RECT -45.490 26.560 94.660 26.700 ;
        RECT 8.010 26.470 8.310 26.560 ;
        RECT 13.760 26.470 14.060 26.560 ;
        RECT 19.510 26.470 19.810 26.560 ;
        RECT 25.260 26.470 25.560 26.560 ;
        RECT 31.010 26.470 31.310 26.560 ;
        RECT 36.760 26.470 37.060 26.560 ;
        RECT 42.510 26.470 42.810 26.560 ;
        RECT 48.260 26.470 48.560 26.560 ;
        RECT 54.010 26.470 54.310 26.560 ;
        RECT 59.760 26.470 60.060 26.560 ;
        RECT 65.510 26.470 65.810 26.560 ;
        RECT 71.260 26.470 71.560 26.560 ;
        RECT 77.010 26.470 77.310 26.560 ;
        RECT 82.760 26.470 83.060 26.560 ;
        RECT 88.510 26.470 88.810 26.560 ;
        RECT 94.260 26.470 94.560 26.560 ;
    END
  END RWLB[4]
  PIN RWL[5]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 25.100 2.760 25.170 ;
        RECT 8.210 25.100 8.510 25.170 ;
        RECT 13.960 25.100 14.260 25.170 ;
        RECT 19.710 25.100 20.010 25.170 ;
        RECT 25.460 25.100 25.760 25.170 ;
        RECT 31.210 25.100 31.510 25.170 ;
        RECT 36.960 25.100 37.260 25.170 ;
        RECT 42.710 25.100 43.010 25.170 ;
        RECT 48.460 25.100 48.760 25.170 ;
        RECT 54.210 25.100 54.510 25.170 ;
        RECT 59.960 25.100 60.260 25.170 ;
        RECT 65.710 25.100 66.010 25.170 ;
        RECT 71.460 25.100 71.760 25.170 ;
        RECT 77.210 25.100 77.510 25.170 ;
        RECT 82.960 25.100 83.260 25.170 ;
        RECT 88.710 25.100 89.010 25.170 ;
        RECT -45.490 24.960 94.660 25.100 ;
        RECT 2.460 24.880 2.760 24.960 ;
        RECT 8.210 24.880 8.510 24.960 ;
        RECT 13.960 24.880 14.260 24.960 ;
        RECT 19.710 24.880 20.010 24.960 ;
        RECT 25.460 24.880 25.760 24.960 ;
        RECT 31.210 24.880 31.510 24.960 ;
        RECT 36.960 24.880 37.260 24.960 ;
        RECT 42.710 24.880 43.010 24.960 ;
        RECT 48.460 24.880 48.760 24.960 ;
        RECT 54.210 24.880 54.510 24.960 ;
        RECT 59.960 24.880 60.260 24.960 ;
        RECT 65.710 24.880 66.010 24.960 ;
        RECT 71.460 24.880 71.760 24.960 ;
        RECT 77.210 24.880 77.510 24.960 ;
        RECT 82.960 24.880 83.260 24.960 ;
        RECT 88.710 24.880 89.010 24.960 ;
    END
  END RWL[5]
  PIN WWL[5]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 24.700 4.730 24.820 ;
        RECT 10.190 24.700 10.480 24.820 ;
        RECT 15.940 24.700 16.230 24.820 ;
        RECT 21.690 24.700 21.980 24.820 ;
        RECT 27.440 24.700 27.730 24.820 ;
        RECT 33.190 24.700 33.480 24.820 ;
        RECT 38.940 24.700 39.230 24.820 ;
        RECT 44.690 24.700 44.980 24.820 ;
        RECT 50.440 24.700 50.730 24.820 ;
        RECT 56.190 24.700 56.480 24.820 ;
        RECT 61.940 24.700 62.230 24.820 ;
        RECT 67.690 24.700 67.980 24.820 ;
        RECT 73.440 24.700 73.730 24.820 ;
        RECT 79.190 24.700 79.480 24.820 ;
        RECT 84.940 24.700 85.230 24.820 ;
        RECT 90.690 24.700 90.980 24.820 ;
        RECT -45.490 24.560 94.660 24.700 ;
        RECT 6.050 24.440 6.340 24.560 ;
        RECT 11.800 24.440 12.090 24.560 ;
        RECT 17.550 24.440 17.840 24.560 ;
        RECT 23.300 24.440 23.590 24.560 ;
        RECT 29.050 24.440 29.340 24.560 ;
        RECT 34.800 24.440 35.090 24.560 ;
        RECT 40.550 24.440 40.840 24.560 ;
        RECT 46.300 24.440 46.590 24.560 ;
        RECT 52.050 24.440 52.340 24.560 ;
        RECT 57.800 24.440 58.090 24.560 ;
        RECT 63.550 24.440 63.840 24.560 ;
        RECT 69.300 24.440 69.590 24.560 ;
        RECT 75.050 24.440 75.340 24.560 ;
        RECT 80.800 24.440 81.090 24.560 ;
        RECT 86.550 24.440 86.840 24.560 ;
        RECT 92.300 24.440 92.590 24.560 ;
    END
  END WWL[5]
  PIN RWLB[5]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 24.290 8.310 24.390 ;
        RECT 13.760 24.290 14.060 24.390 ;
        RECT 19.510 24.290 19.810 24.390 ;
        RECT 25.260 24.290 25.560 24.390 ;
        RECT 31.010 24.290 31.310 24.390 ;
        RECT 36.760 24.290 37.060 24.390 ;
        RECT 42.510 24.290 42.810 24.390 ;
        RECT 48.260 24.290 48.560 24.390 ;
        RECT 54.010 24.290 54.310 24.390 ;
        RECT 59.760 24.290 60.060 24.390 ;
        RECT 65.510 24.290 65.810 24.390 ;
        RECT 71.260 24.290 71.560 24.390 ;
        RECT 77.010 24.290 77.310 24.390 ;
        RECT 82.760 24.290 83.060 24.390 ;
        RECT 88.510 24.290 88.810 24.390 ;
        RECT 94.260 24.290 94.560 24.390 ;
        RECT -45.490 24.150 94.660 24.290 ;
        RECT 8.010 24.060 8.310 24.150 ;
        RECT 13.760 24.060 14.060 24.150 ;
        RECT 19.510 24.060 19.810 24.150 ;
        RECT 25.260 24.060 25.560 24.150 ;
        RECT 31.010 24.060 31.310 24.150 ;
        RECT 36.760 24.060 37.060 24.150 ;
        RECT 42.510 24.060 42.810 24.150 ;
        RECT 48.260 24.060 48.560 24.150 ;
        RECT 54.010 24.060 54.310 24.150 ;
        RECT 59.760 24.060 60.060 24.150 ;
        RECT 65.510 24.060 65.810 24.150 ;
        RECT 71.260 24.060 71.560 24.150 ;
        RECT 77.010 24.060 77.310 24.150 ;
        RECT 82.760 24.060 83.060 24.150 ;
        RECT 88.510 24.060 88.810 24.150 ;
        RECT 94.260 24.060 94.560 24.150 ;
    END
  END RWLB[5]
  PIN RWL[6]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 22.690 2.760 22.760 ;
        RECT 8.210 22.690 8.510 22.760 ;
        RECT 13.960 22.690 14.260 22.760 ;
        RECT 19.710 22.690 20.010 22.760 ;
        RECT 25.460 22.690 25.760 22.760 ;
        RECT 31.210 22.690 31.510 22.760 ;
        RECT 36.960 22.690 37.260 22.760 ;
        RECT 42.710 22.690 43.010 22.760 ;
        RECT 48.460 22.690 48.760 22.760 ;
        RECT 54.210 22.690 54.510 22.760 ;
        RECT 59.960 22.690 60.260 22.760 ;
        RECT 65.710 22.690 66.010 22.760 ;
        RECT 71.460 22.690 71.760 22.760 ;
        RECT 77.210 22.690 77.510 22.760 ;
        RECT 82.960 22.690 83.260 22.760 ;
        RECT 88.710 22.690 89.010 22.760 ;
        RECT -45.490 22.550 94.660 22.690 ;
        RECT 2.460 22.470 2.760 22.550 ;
        RECT 8.210 22.470 8.510 22.550 ;
        RECT 13.960 22.470 14.260 22.550 ;
        RECT 19.710 22.470 20.010 22.550 ;
        RECT 25.460 22.470 25.760 22.550 ;
        RECT 31.210 22.470 31.510 22.550 ;
        RECT 36.960 22.470 37.260 22.550 ;
        RECT 42.710 22.470 43.010 22.550 ;
        RECT 48.460 22.470 48.760 22.550 ;
        RECT 54.210 22.470 54.510 22.550 ;
        RECT 59.960 22.470 60.260 22.550 ;
        RECT 65.710 22.470 66.010 22.550 ;
        RECT 71.460 22.470 71.760 22.550 ;
        RECT 77.210 22.470 77.510 22.550 ;
        RECT 82.960 22.470 83.260 22.550 ;
        RECT 88.710 22.470 89.010 22.550 ;
    END
  END RWL[6]
  PIN WWL[6]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 22.290 4.730 22.410 ;
        RECT 10.190 22.290 10.480 22.410 ;
        RECT 15.940 22.290 16.230 22.410 ;
        RECT 21.690 22.290 21.980 22.410 ;
        RECT 27.440 22.290 27.730 22.410 ;
        RECT 33.190 22.290 33.480 22.410 ;
        RECT 38.940 22.290 39.230 22.410 ;
        RECT 44.690 22.290 44.980 22.410 ;
        RECT 50.440 22.290 50.730 22.410 ;
        RECT 56.190 22.290 56.480 22.410 ;
        RECT 61.940 22.290 62.230 22.410 ;
        RECT 67.690 22.290 67.980 22.410 ;
        RECT 73.440 22.290 73.730 22.410 ;
        RECT 79.190 22.290 79.480 22.410 ;
        RECT 84.940 22.290 85.230 22.410 ;
        RECT 90.690 22.290 90.980 22.410 ;
        RECT -45.490 22.150 94.660 22.290 ;
        RECT 6.050 22.030 6.340 22.150 ;
        RECT 11.800 22.030 12.090 22.150 ;
        RECT 17.550 22.030 17.840 22.150 ;
        RECT 23.300 22.030 23.590 22.150 ;
        RECT 29.050 22.030 29.340 22.150 ;
        RECT 34.800 22.030 35.090 22.150 ;
        RECT 40.550 22.030 40.840 22.150 ;
        RECT 46.300 22.030 46.590 22.150 ;
        RECT 52.050 22.030 52.340 22.150 ;
        RECT 57.800 22.030 58.090 22.150 ;
        RECT 63.550 22.030 63.840 22.150 ;
        RECT 69.300 22.030 69.590 22.150 ;
        RECT 75.050 22.030 75.340 22.150 ;
        RECT 80.800 22.030 81.090 22.150 ;
        RECT 86.550 22.030 86.840 22.150 ;
        RECT 92.300 22.030 92.590 22.150 ;
    END
  END WWL[6]
  PIN RWLB[6]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 21.880 8.310 21.980 ;
        RECT 13.760 21.880 14.060 21.980 ;
        RECT 19.510 21.880 19.810 21.980 ;
        RECT 25.260 21.880 25.560 21.980 ;
        RECT 31.010 21.880 31.310 21.980 ;
        RECT 36.760 21.880 37.060 21.980 ;
        RECT 42.510 21.880 42.810 21.980 ;
        RECT 48.260 21.880 48.560 21.980 ;
        RECT 54.010 21.880 54.310 21.980 ;
        RECT 59.760 21.880 60.060 21.980 ;
        RECT 65.510 21.880 65.810 21.980 ;
        RECT 71.260 21.880 71.560 21.980 ;
        RECT 77.010 21.880 77.310 21.980 ;
        RECT 82.760 21.880 83.060 21.980 ;
        RECT 88.510 21.880 88.810 21.980 ;
        RECT 94.260 21.880 94.560 21.980 ;
        RECT -45.490 21.740 94.660 21.880 ;
        RECT 8.010 21.650 8.310 21.740 ;
        RECT 13.760 21.650 14.060 21.740 ;
        RECT 19.510 21.650 19.810 21.740 ;
        RECT 25.260 21.650 25.560 21.740 ;
        RECT 31.010 21.650 31.310 21.740 ;
        RECT 36.760 21.650 37.060 21.740 ;
        RECT 42.510 21.650 42.810 21.740 ;
        RECT 48.260 21.650 48.560 21.740 ;
        RECT 54.010 21.650 54.310 21.740 ;
        RECT 59.760 21.650 60.060 21.740 ;
        RECT 65.510 21.650 65.810 21.740 ;
        RECT 71.260 21.650 71.560 21.740 ;
        RECT 77.010 21.650 77.310 21.740 ;
        RECT 82.760 21.650 83.060 21.740 ;
        RECT 88.510 21.650 88.810 21.740 ;
        RECT 94.260 21.650 94.560 21.740 ;
    END
  END RWLB[6]
  PIN RWL[7]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 20.280 2.760 20.350 ;
        RECT 8.210 20.280 8.510 20.350 ;
        RECT 13.960 20.280 14.260 20.350 ;
        RECT 19.710 20.280 20.010 20.350 ;
        RECT 25.460 20.280 25.760 20.350 ;
        RECT 31.210 20.280 31.510 20.350 ;
        RECT 36.960 20.280 37.260 20.350 ;
        RECT 42.710 20.280 43.010 20.350 ;
        RECT 48.460 20.280 48.760 20.350 ;
        RECT 54.210 20.280 54.510 20.350 ;
        RECT 59.960 20.280 60.260 20.350 ;
        RECT 65.710 20.280 66.010 20.350 ;
        RECT 71.460 20.280 71.760 20.350 ;
        RECT 77.210 20.280 77.510 20.350 ;
        RECT 82.960 20.280 83.260 20.350 ;
        RECT 88.710 20.280 89.010 20.350 ;
        RECT -45.490 20.140 94.660 20.280 ;
        RECT 2.460 20.060 2.760 20.140 ;
        RECT 8.210 20.060 8.510 20.140 ;
        RECT 13.960 20.060 14.260 20.140 ;
        RECT 19.710 20.060 20.010 20.140 ;
        RECT 25.460 20.060 25.760 20.140 ;
        RECT 31.210 20.060 31.510 20.140 ;
        RECT 36.960 20.060 37.260 20.140 ;
        RECT 42.710 20.060 43.010 20.140 ;
        RECT 48.460 20.060 48.760 20.140 ;
        RECT 54.210 20.060 54.510 20.140 ;
        RECT 59.960 20.060 60.260 20.140 ;
        RECT 65.710 20.060 66.010 20.140 ;
        RECT 71.460 20.060 71.760 20.140 ;
        RECT 77.210 20.060 77.510 20.140 ;
        RECT 82.960 20.060 83.260 20.140 ;
        RECT 88.710 20.060 89.010 20.140 ;
    END
  END RWL[7]
  PIN WWL[7]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 19.880 4.730 20.000 ;
        RECT 10.190 19.880 10.480 20.000 ;
        RECT 15.940 19.880 16.230 20.000 ;
        RECT 21.690 19.880 21.980 20.000 ;
        RECT 27.440 19.880 27.730 20.000 ;
        RECT 33.190 19.880 33.480 20.000 ;
        RECT 38.940 19.880 39.230 20.000 ;
        RECT 44.690 19.880 44.980 20.000 ;
        RECT 50.440 19.880 50.730 20.000 ;
        RECT 56.190 19.880 56.480 20.000 ;
        RECT 61.940 19.880 62.230 20.000 ;
        RECT 67.690 19.880 67.980 20.000 ;
        RECT 73.440 19.880 73.730 20.000 ;
        RECT 79.190 19.880 79.480 20.000 ;
        RECT 84.940 19.880 85.230 20.000 ;
        RECT 90.690 19.880 90.980 20.000 ;
        RECT -45.490 19.740 94.660 19.880 ;
        RECT 6.050 19.620 6.340 19.740 ;
        RECT 11.800 19.620 12.090 19.740 ;
        RECT 17.550 19.620 17.840 19.740 ;
        RECT 23.300 19.620 23.590 19.740 ;
        RECT 29.050 19.620 29.340 19.740 ;
        RECT 34.800 19.620 35.090 19.740 ;
        RECT 40.550 19.620 40.840 19.740 ;
        RECT 46.300 19.620 46.590 19.740 ;
        RECT 52.050 19.620 52.340 19.740 ;
        RECT 57.800 19.620 58.090 19.740 ;
        RECT 63.550 19.620 63.840 19.740 ;
        RECT 69.300 19.620 69.590 19.740 ;
        RECT 75.050 19.620 75.340 19.740 ;
        RECT 80.800 19.620 81.090 19.740 ;
        RECT 86.550 19.620 86.840 19.740 ;
        RECT 92.300 19.620 92.590 19.740 ;
    END
  END WWL[7]
  PIN RWLB[7]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 19.470 8.310 19.570 ;
        RECT 13.760 19.470 14.060 19.570 ;
        RECT 19.510 19.470 19.810 19.570 ;
        RECT 25.260 19.470 25.560 19.570 ;
        RECT 31.010 19.470 31.310 19.570 ;
        RECT 36.760 19.470 37.060 19.570 ;
        RECT 42.510 19.470 42.810 19.570 ;
        RECT 48.260 19.470 48.560 19.570 ;
        RECT 54.010 19.470 54.310 19.570 ;
        RECT 59.760 19.470 60.060 19.570 ;
        RECT 65.510 19.470 65.810 19.570 ;
        RECT 71.260 19.470 71.560 19.570 ;
        RECT 77.010 19.470 77.310 19.570 ;
        RECT 82.760 19.470 83.060 19.570 ;
        RECT 88.510 19.470 88.810 19.570 ;
        RECT 94.260 19.470 94.560 19.570 ;
        RECT -45.490 19.330 94.660 19.470 ;
        RECT 8.010 19.240 8.310 19.330 ;
        RECT 13.760 19.240 14.060 19.330 ;
        RECT 19.510 19.240 19.810 19.330 ;
        RECT 25.260 19.240 25.560 19.330 ;
        RECT 31.010 19.240 31.310 19.330 ;
        RECT 36.760 19.240 37.060 19.330 ;
        RECT 42.510 19.240 42.810 19.330 ;
        RECT 48.260 19.240 48.560 19.330 ;
        RECT 54.010 19.240 54.310 19.330 ;
        RECT 59.760 19.240 60.060 19.330 ;
        RECT 65.510 19.240 65.810 19.330 ;
        RECT 71.260 19.240 71.560 19.330 ;
        RECT 77.010 19.240 77.310 19.330 ;
        RECT 82.760 19.240 83.060 19.330 ;
        RECT 88.510 19.240 88.810 19.330 ;
        RECT 94.260 19.240 94.560 19.330 ;
    END
  END RWLB[7]
  PIN RWL[8]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 17.870 2.760 17.940 ;
        RECT 8.210 17.870 8.510 17.940 ;
        RECT 13.960 17.870 14.260 17.940 ;
        RECT 19.710 17.870 20.010 17.940 ;
        RECT 25.460 17.870 25.760 17.940 ;
        RECT 31.210 17.870 31.510 17.940 ;
        RECT 36.960 17.870 37.260 17.940 ;
        RECT 42.710 17.870 43.010 17.940 ;
        RECT 48.460 17.870 48.760 17.940 ;
        RECT 54.210 17.870 54.510 17.940 ;
        RECT 59.960 17.870 60.260 17.940 ;
        RECT 65.710 17.870 66.010 17.940 ;
        RECT 71.460 17.870 71.760 17.940 ;
        RECT 77.210 17.870 77.510 17.940 ;
        RECT 82.960 17.870 83.260 17.940 ;
        RECT 88.710 17.870 89.010 17.940 ;
        RECT -45.490 17.730 94.660 17.870 ;
        RECT 2.460 17.650 2.760 17.730 ;
        RECT 8.210 17.650 8.510 17.730 ;
        RECT 13.960 17.650 14.260 17.730 ;
        RECT 19.710 17.650 20.010 17.730 ;
        RECT 25.460 17.650 25.760 17.730 ;
        RECT 31.210 17.650 31.510 17.730 ;
        RECT 36.960 17.650 37.260 17.730 ;
        RECT 42.710 17.650 43.010 17.730 ;
        RECT 48.460 17.650 48.760 17.730 ;
        RECT 54.210 17.650 54.510 17.730 ;
        RECT 59.960 17.650 60.260 17.730 ;
        RECT 65.710 17.650 66.010 17.730 ;
        RECT 71.460 17.650 71.760 17.730 ;
        RECT 77.210 17.650 77.510 17.730 ;
        RECT 82.960 17.650 83.260 17.730 ;
        RECT 88.710 17.650 89.010 17.730 ;
    END
  END RWL[8]
  PIN WWL[8]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 17.470 4.730 17.590 ;
        RECT 10.190 17.470 10.480 17.590 ;
        RECT 15.940 17.470 16.230 17.590 ;
        RECT 21.690 17.470 21.980 17.590 ;
        RECT 27.440 17.470 27.730 17.590 ;
        RECT 33.190 17.470 33.480 17.590 ;
        RECT 38.940 17.470 39.230 17.590 ;
        RECT 44.690 17.470 44.980 17.590 ;
        RECT 50.440 17.470 50.730 17.590 ;
        RECT 56.190 17.470 56.480 17.590 ;
        RECT 61.940 17.470 62.230 17.590 ;
        RECT 67.690 17.470 67.980 17.590 ;
        RECT 73.440 17.470 73.730 17.590 ;
        RECT 79.190 17.470 79.480 17.590 ;
        RECT 84.940 17.470 85.230 17.590 ;
        RECT 90.690 17.470 90.980 17.590 ;
        RECT -45.490 17.330 94.660 17.470 ;
        RECT 6.050 17.210 6.340 17.330 ;
        RECT 11.800 17.210 12.090 17.330 ;
        RECT 17.550 17.210 17.840 17.330 ;
        RECT 23.300 17.210 23.590 17.330 ;
        RECT 29.050 17.210 29.340 17.330 ;
        RECT 34.800 17.210 35.090 17.330 ;
        RECT 40.550 17.210 40.840 17.330 ;
        RECT 46.300 17.210 46.590 17.330 ;
        RECT 52.050 17.210 52.340 17.330 ;
        RECT 57.800 17.210 58.090 17.330 ;
        RECT 63.550 17.210 63.840 17.330 ;
        RECT 69.300 17.210 69.590 17.330 ;
        RECT 75.050 17.210 75.340 17.330 ;
        RECT 80.800 17.210 81.090 17.330 ;
        RECT 86.550 17.210 86.840 17.330 ;
        RECT 92.300 17.210 92.590 17.330 ;
    END
  END WWL[8]
  PIN RWLB[8]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 17.060 8.310 17.160 ;
        RECT 13.760 17.060 14.060 17.160 ;
        RECT 19.510 17.060 19.810 17.160 ;
        RECT 25.260 17.060 25.560 17.160 ;
        RECT 31.010 17.060 31.310 17.160 ;
        RECT 36.760 17.060 37.060 17.160 ;
        RECT 42.510 17.060 42.810 17.160 ;
        RECT 48.260 17.060 48.560 17.160 ;
        RECT 54.010 17.060 54.310 17.160 ;
        RECT 59.760 17.060 60.060 17.160 ;
        RECT 65.510 17.060 65.810 17.160 ;
        RECT 71.260 17.060 71.560 17.160 ;
        RECT 77.010 17.060 77.310 17.160 ;
        RECT 82.760 17.060 83.060 17.160 ;
        RECT 88.510 17.060 88.810 17.160 ;
        RECT 94.260 17.060 94.560 17.160 ;
        RECT -45.490 16.920 94.660 17.060 ;
        RECT 8.010 16.830 8.310 16.920 ;
        RECT 13.760 16.830 14.060 16.920 ;
        RECT 19.510 16.830 19.810 16.920 ;
        RECT 25.260 16.830 25.560 16.920 ;
        RECT 31.010 16.830 31.310 16.920 ;
        RECT 36.760 16.830 37.060 16.920 ;
        RECT 42.510 16.830 42.810 16.920 ;
        RECT 48.260 16.830 48.560 16.920 ;
        RECT 54.010 16.830 54.310 16.920 ;
        RECT 59.760 16.830 60.060 16.920 ;
        RECT 65.510 16.830 65.810 16.920 ;
        RECT 71.260 16.830 71.560 16.920 ;
        RECT 77.010 16.830 77.310 16.920 ;
        RECT 82.760 16.830 83.060 16.920 ;
        RECT 88.510 16.830 88.810 16.920 ;
        RECT 94.260 16.830 94.560 16.920 ;
    END
  END RWLB[8]
  PIN RWL[9]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 15.460 2.760 15.530 ;
        RECT 8.210 15.460 8.510 15.530 ;
        RECT 13.960 15.460 14.260 15.530 ;
        RECT 19.710 15.460 20.010 15.530 ;
        RECT 25.460 15.460 25.760 15.530 ;
        RECT 31.210 15.460 31.510 15.530 ;
        RECT 36.960 15.460 37.260 15.530 ;
        RECT 42.710 15.460 43.010 15.530 ;
        RECT 48.460 15.460 48.760 15.530 ;
        RECT 54.210 15.460 54.510 15.530 ;
        RECT 59.960 15.460 60.260 15.530 ;
        RECT 65.710 15.460 66.010 15.530 ;
        RECT 71.460 15.460 71.760 15.530 ;
        RECT 77.210 15.460 77.510 15.530 ;
        RECT 82.960 15.460 83.260 15.530 ;
        RECT 88.710 15.460 89.010 15.530 ;
        RECT -45.490 15.320 94.660 15.460 ;
        RECT 2.460 15.240 2.760 15.320 ;
        RECT 8.210 15.240 8.510 15.320 ;
        RECT 13.960 15.240 14.260 15.320 ;
        RECT 19.710 15.240 20.010 15.320 ;
        RECT 25.460 15.240 25.760 15.320 ;
        RECT 31.210 15.240 31.510 15.320 ;
        RECT 36.960 15.240 37.260 15.320 ;
        RECT 42.710 15.240 43.010 15.320 ;
        RECT 48.460 15.240 48.760 15.320 ;
        RECT 54.210 15.240 54.510 15.320 ;
        RECT 59.960 15.240 60.260 15.320 ;
        RECT 65.710 15.240 66.010 15.320 ;
        RECT 71.460 15.240 71.760 15.320 ;
        RECT 77.210 15.240 77.510 15.320 ;
        RECT 82.960 15.240 83.260 15.320 ;
        RECT 88.710 15.240 89.010 15.320 ;
    END
  END RWL[9]
  PIN WWL[9]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 15.060 4.730 15.180 ;
        RECT 10.190 15.060 10.480 15.180 ;
        RECT 15.940 15.060 16.230 15.180 ;
        RECT 21.690 15.060 21.980 15.180 ;
        RECT 27.440 15.060 27.730 15.180 ;
        RECT 33.190 15.060 33.480 15.180 ;
        RECT 38.940 15.060 39.230 15.180 ;
        RECT 44.690 15.060 44.980 15.180 ;
        RECT 50.440 15.060 50.730 15.180 ;
        RECT 56.190 15.060 56.480 15.180 ;
        RECT 61.940 15.060 62.230 15.180 ;
        RECT 67.690 15.060 67.980 15.180 ;
        RECT 73.440 15.060 73.730 15.180 ;
        RECT 79.190 15.060 79.480 15.180 ;
        RECT 84.940 15.060 85.230 15.180 ;
        RECT 90.690 15.060 90.980 15.180 ;
        RECT -45.490 14.920 94.660 15.060 ;
        RECT 6.050 14.800 6.340 14.920 ;
        RECT 11.800 14.800 12.090 14.920 ;
        RECT 17.550 14.800 17.840 14.920 ;
        RECT 23.300 14.800 23.590 14.920 ;
        RECT 29.050 14.800 29.340 14.920 ;
        RECT 34.800 14.800 35.090 14.920 ;
        RECT 40.550 14.800 40.840 14.920 ;
        RECT 46.300 14.800 46.590 14.920 ;
        RECT 52.050 14.800 52.340 14.920 ;
        RECT 57.800 14.800 58.090 14.920 ;
        RECT 63.550 14.800 63.840 14.920 ;
        RECT 69.300 14.800 69.590 14.920 ;
        RECT 75.050 14.800 75.340 14.920 ;
        RECT 80.800 14.800 81.090 14.920 ;
        RECT 86.550 14.800 86.840 14.920 ;
        RECT 92.300 14.800 92.590 14.920 ;
    END
  END WWL[9]
  PIN RWLB[9]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 14.650 8.310 14.750 ;
        RECT 13.760 14.650 14.060 14.750 ;
        RECT 19.510 14.650 19.810 14.750 ;
        RECT 25.260 14.650 25.560 14.750 ;
        RECT 31.010 14.650 31.310 14.750 ;
        RECT 36.760 14.650 37.060 14.750 ;
        RECT 42.510 14.650 42.810 14.750 ;
        RECT 48.260 14.650 48.560 14.750 ;
        RECT 54.010 14.650 54.310 14.750 ;
        RECT 59.760 14.650 60.060 14.750 ;
        RECT 65.510 14.650 65.810 14.750 ;
        RECT 71.260 14.650 71.560 14.750 ;
        RECT 77.010 14.650 77.310 14.750 ;
        RECT 82.760 14.650 83.060 14.750 ;
        RECT 88.510 14.650 88.810 14.750 ;
        RECT 94.260 14.650 94.560 14.750 ;
        RECT -45.490 14.510 94.660 14.650 ;
        RECT 8.010 14.420 8.310 14.510 ;
        RECT 13.760 14.420 14.060 14.510 ;
        RECT 19.510 14.420 19.810 14.510 ;
        RECT 25.260 14.420 25.560 14.510 ;
        RECT 31.010 14.420 31.310 14.510 ;
        RECT 36.760 14.420 37.060 14.510 ;
        RECT 42.510 14.420 42.810 14.510 ;
        RECT 48.260 14.420 48.560 14.510 ;
        RECT 54.010 14.420 54.310 14.510 ;
        RECT 59.760 14.420 60.060 14.510 ;
        RECT 65.510 14.420 65.810 14.510 ;
        RECT 71.260 14.420 71.560 14.510 ;
        RECT 77.010 14.420 77.310 14.510 ;
        RECT 82.760 14.420 83.060 14.510 ;
        RECT 88.510 14.420 88.810 14.510 ;
        RECT 94.260 14.420 94.560 14.510 ;
    END
  END RWLB[9]
  PIN RWL[10]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 13.050 2.760 13.120 ;
        RECT 8.210 13.050 8.510 13.120 ;
        RECT 13.960 13.050 14.260 13.120 ;
        RECT 19.710 13.050 20.010 13.120 ;
        RECT 25.460 13.050 25.760 13.120 ;
        RECT 31.210 13.050 31.510 13.120 ;
        RECT 36.960 13.050 37.260 13.120 ;
        RECT 42.710 13.050 43.010 13.120 ;
        RECT 48.460 13.050 48.760 13.120 ;
        RECT 54.210 13.050 54.510 13.120 ;
        RECT 59.960 13.050 60.260 13.120 ;
        RECT 65.710 13.050 66.010 13.120 ;
        RECT 71.460 13.050 71.760 13.120 ;
        RECT 77.210 13.050 77.510 13.120 ;
        RECT 82.960 13.050 83.260 13.120 ;
        RECT 88.710 13.050 89.010 13.120 ;
        RECT -45.490 12.910 94.660 13.050 ;
        RECT 2.460 12.830 2.760 12.910 ;
        RECT 8.210 12.830 8.510 12.910 ;
        RECT 13.960 12.830 14.260 12.910 ;
        RECT 19.710 12.830 20.010 12.910 ;
        RECT 25.460 12.830 25.760 12.910 ;
        RECT 31.210 12.830 31.510 12.910 ;
        RECT 36.960 12.830 37.260 12.910 ;
        RECT 42.710 12.830 43.010 12.910 ;
        RECT 48.460 12.830 48.760 12.910 ;
        RECT 54.210 12.830 54.510 12.910 ;
        RECT 59.960 12.830 60.260 12.910 ;
        RECT 65.710 12.830 66.010 12.910 ;
        RECT 71.460 12.830 71.760 12.910 ;
        RECT 77.210 12.830 77.510 12.910 ;
        RECT 82.960 12.830 83.260 12.910 ;
        RECT 88.710 12.830 89.010 12.910 ;
    END
  END RWL[10]
  PIN WWL[10]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 12.650 4.730 12.770 ;
        RECT 10.190 12.650 10.480 12.770 ;
        RECT 15.940 12.650 16.230 12.770 ;
        RECT 21.690 12.650 21.980 12.770 ;
        RECT 27.440 12.650 27.730 12.770 ;
        RECT 33.190 12.650 33.480 12.770 ;
        RECT 38.940 12.650 39.230 12.770 ;
        RECT 44.690 12.650 44.980 12.770 ;
        RECT 50.440 12.650 50.730 12.770 ;
        RECT 56.190 12.650 56.480 12.770 ;
        RECT 61.940 12.650 62.230 12.770 ;
        RECT 67.690 12.650 67.980 12.770 ;
        RECT 73.440 12.650 73.730 12.770 ;
        RECT 79.190 12.650 79.480 12.770 ;
        RECT 84.940 12.650 85.230 12.770 ;
        RECT 90.690 12.650 90.980 12.770 ;
        RECT -45.490 12.510 94.660 12.650 ;
        RECT 6.050 12.390 6.340 12.510 ;
        RECT 11.800 12.390 12.090 12.510 ;
        RECT 17.550 12.390 17.840 12.510 ;
        RECT 23.300 12.390 23.590 12.510 ;
        RECT 29.050 12.390 29.340 12.510 ;
        RECT 34.800 12.390 35.090 12.510 ;
        RECT 40.550 12.390 40.840 12.510 ;
        RECT 46.300 12.390 46.590 12.510 ;
        RECT 52.050 12.390 52.340 12.510 ;
        RECT 57.800 12.390 58.090 12.510 ;
        RECT 63.550 12.390 63.840 12.510 ;
        RECT 69.300 12.390 69.590 12.510 ;
        RECT 75.050 12.390 75.340 12.510 ;
        RECT 80.800 12.390 81.090 12.510 ;
        RECT 86.550 12.390 86.840 12.510 ;
        RECT 92.300 12.390 92.590 12.510 ;
    END
  END WWL[10]
  PIN RWLB[10]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 12.240 8.310 12.340 ;
        RECT 13.760 12.240 14.060 12.340 ;
        RECT 19.510 12.240 19.810 12.340 ;
        RECT 25.260 12.240 25.560 12.340 ;
        RECT 31.010 12.240 31.310 12.340 ;
        RECT 36.760 12.240 37.060 12.340 ;
        RECT 42.510 12.240 42.810 12.340 ;
        RECT 48.260 12.240 48.560 12.340 ;
        RECT 54.010 12.240 54.310 12.340 ;
        RECT 59.760 12.240 60.060 12.340 ;
        RECT 65.510 12.240 65.810 12.340 ;
        RECT 71.260 12.240 71.560 12.340 ;
        RECT 77.010 12.240 77.310 12.340 ;
        RECT 82.760 12.240 83.060 12.340 ;
        RECT 88.510 12.240 88.810 12.340 ;
        RECT 94.260 12.240 94.560 12.340 ;
        RECT -45.490 12.100 94.660 12.240 ;
        RECT 8.010 12.010 8.310 12.100 ;
        RECT 13.760 12.010 14.060 12.100 ;
        RECT 19.510 12.010 19.810 12.100 ;
        RECT 25.260 12.010 25.560 12.100 ;
        RECT 31.010 12.010 31.310 12.100 ;
        RECT 36.760 12.010 37.060 12.100 ;
        RECT 42.510 12.010 42.810 12.100 ;
        RECT 48.260 12.010 48.560 12.100 ;
        RECT 54.010 12.010 54.310 12.100 ;
        RECT 59.760 12.010 60.060 12.100 ;
        RECT 65.510 12.010 65.810 12.100 ;
        RECT 71.260 12.010 71.560 12.100 ;
        RECT 77.010 12.010 77.310 12.100 ;
        RECT 82.760 12.010 83.060 12.100 ;
        RECT 88.510 12.010 88.810 12.100 ;
        RECT 94.260 12.010 94.560 12.100 ;
    END
  END RWLB[10]
  PIN RWL[11]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 10.640 2.760 10.710 ;
        RECT 8.210 10.640 8.510 10.710 ;
        RECT 13.960 10.640 14.260 10.710 ;
        RECT 19.710 10.640 20.010 10.710 ;
        RECT 25.460 10.640 25.760 10.710 ;
        RECT 31.210 10.640 31.510 10.710 ;
        RECT 36.960 10.640 37.260 10.710 ;
        RECT 42.710 10.640 43.010 10.710 ;
        RECT 48.460 10.640 48.760 10.710 ;
        RECT 54.210 10.640 54.510 10.710 ;
        RECT 59.960 10.640 60.260 10.710 ;
        RECT 65.710 10.640 66.010 10.710 ;
        RECT 71.460 10.640 71.760 10.710 ;
        RECT 77.210 10.640 77.510 10.710 ;
        RECT 82.960 10.640 83.260 10.710 ;
        RECT 88.710 10.640 89.010 10.710 ;
        RECT -45.490 10.500 94.660 10.640 ;
        RECT 2.460 10.420 2.760 10.500 ;
        RECT 8.210 10.420 8.510 10.500 ;
        RECT 13.960 10.420 14.260 10.500 ;
        RECT 19.710 10.420 20.010 10.500 ;
        RECT 25.460 10.420 25.760 10.500 ;
        RECT 31.210 10.420 31.510 10.500 ;
        RECT 36.960 10.420 37.260 10.500 ;
        RECT 42.710 10.420 43.010 10.500 ;
        RECT 48.460 10.420 48.760 10.500 ;
        RECT 54.210 10.420 54.510 10.500 ;
        RECT 59.960 10.420 60.260 10.500 ;
        RECT 65.710 10.420 66.010 10.500 ;
        RECT 71.460 10.420 71.760 10.500 ;
        RECT 77.210 10.420 77.510 10.500 ;
        RECT 82.960 10.420 83.260 10.500 ;
        RECT 88.710 10.420 89.010 10.500 ;
    END
  END RWL[11]
  PIN WWL[11]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 10.240 4.730 10.360 ;
        RECT 10.190 10.240 10.480 10.360 ;
        RECT 15.940 10.240 16.230 10.360 ;
        RECT 21.690 10.240 21.980 10.360 ;
        RECT 27.440 10.240 27.730 10.360 ;
        RECT 33.190 10.240 33.480 10.360 ;
        RECT 38.940 10.240 39.230 10.360 ;
        RECT 44.690 10.240 44.980 10.360 ;
        RECT 50.440 10.240 50.730 10.360 ;
        RECT 56.190 10.240 56.480 10.360 ;
        RECT 61.940 10.240 62.230 10.360 ;
        RECT 67.690 10.240 67.980 10.360 ;
        RECT 73.440 10.240 73.730 10.360 ;
        RECT 79.190 10.240 79.480 10.360 ;
        RECT 84.940 10.240 85.230 10.360 ;
        RECT 90.690 10.240 90.980 10.360 ;
        RECT -45.490 10.100 94.660 10.240 ;
        RECT 6.050 9.980 6.340 10.100 ;
        RECT 11.800 9.980 12.090 10.100 ;
        RECT 17.550 9.980 17.840 10.100 ;
        RECT 23.300 9.980 23.590 10.100 ;
        RECT 29.050 9.980 29.340 10.100 ;
        RECT 34.800 9.980 35.090 10.100 ;
        RECT 40.550 9.980 40.840 10.100 ;
        RECT 46.300 9.980 46.590 10.100 ;
        RECT 52.050 9.980 52.340 10.100 ;
        RECT 57.800 9.980 58.090 10.100 ;
        RECT 63.550 9.980 63.840 10.100 ;
        RECT 69.300 9.980 69.590 10.100 ;
        RECT 75.050 9.980 75.340 10.100 ;
        RECT 80.800 9.980 81.090 10.100 ;
        RECT 86.550 9.980 86.840 10.100 ;
        RECT 92.300 9.980 92.590 10.100 ;
    END
  END WWL[11]
  PIN RWLB[11]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 9.830 8.310 9.930 ;
        RECT 13.760 9.830 14.060 9.930 ;
        RECT 19.510 9.830 19.810 9.930 ;
        RECT 25.260 9.830 25.560 9.930 ;
        RECT 31.010 9.830 31.310 9.930 ;
        RECT 36.760 9.830 37.060 9.930 ;
        RECT 42.510 9.830 42.810 9.930 ;
        RECT 48.260 9.830 48.560 9.930 ;
        RECT 54.010 9.830 54.310 9.930 ;
        RECT 59.760 9.830 60.060 9.930 ;
        RECT 65.510 9.830 65.810 9.930 ;
        RECT 71.260 9.830 71.560 9.930 ;
        RECT 77.010 9.830 77.310 9.930 ;
        RECT 82.760 9.830 83.060 9.930 ;
        RECT 88.510 9.830 88.810 9.930 ;
        RECT 94.260 9.830 94.560 9.930 ;
        RECT -45.490 9.690 94.660 9.830 ;
        RECT 8.010 9.600 8.310 9.690 ;
        RECT 13.760 9.600 14.060 9.690 ;
        RECT 19.510 9.600 19.810 9.690 ;
        RECT 25.260 9.600 25.560 9.690 ;
        RECT 31.010 9.600 31.310 9.690 ;
        RECT 36.760 9.600 37.060 9.690 ;
        RECT 42.510 9.600 42.810 9.690 ;
        RECT 48.260 9.600 48.560 9.690 ;
        RECT 54.010 9.600 54.310 9.690 ;
        RECT 59.760 9.600 60.060 9.690 ;
        RECT 65.510 9.600 65.810 9.690 ;
        RECT 71.260 9.600 71.560 9.690 ;
        RECT 77.010 9.600 77.310 9.690 ;
        RECT 82.760 9.600 83.060 9.690 ;
        RECT 88.510 9.600 88.810 9.690 ;
        RECT 94.260 9.600 94.560 9.690 ;
    END
  END RWLB[11]
  PIN RWL[12]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 7.820 2.760 7.880 ;
        RECT 8.210 7.820 8.510 7.880 ;
        RECT 13.960 7.820 14.260 7.880 ;
        RECT 19.710 7.820 20.010 7.880 ;
        RECT 25.460 7.820 25.760 7.880 ;
        RECT 31.210 7.820 31.510 7.880 ;
        RECT 36.960 7.820 37.260 7.880 ;
        RECT 42.710 7.820 43.010 7.880 ;
        RECT 48.460 7.820 48.760 7.880 ;
        RECT 54.210 7.820 54.510 7.880 ;
        RECT 59.960 7.820 60.260 7.880 ;
        RECT 65.710 7.820 66.010 7.880 ;
        RECT 71.460 7.820 71.760 7.880 ;
        RECT 77.210 7.820 77.510 7.880 ;
        RECT 82.960 7.820 83.260 7.880 ;
        RECT 88.710 7.820 89.010 7.880 ;
        RECT -45.490 7.680 94.660 7.820 ;
        RECT 2.460 7.600 2.760 7.680 ;
        RECT 8.210 7.600 8.510 7.680 ;
        RECT 13.960 7.600 14.260 7.680 ;
        RECT 19.710 7.600 20.010 7.680 ;
        RECT 25.460 7.600 25.760 7.680 ;
        RECT 31.210 7.600 31.510 7.680 ;
        RECT 36.960 7.600 37.260 7.680 ;
        RECT 42.710 7.600 43.010 7.680 ;
        RECT 48.460 7.600 48.760 7.680 ;
        RECT 54.210 7.600 54.510 7.680 ;
        RECT 59.960 7.600 60.260 7.680 ;
        RECT 65.710 7.600 66.010 7.680 ;
        RECT 71.460 7.600 71.760 7.680 ;
        RECT 77.210 7.600 77.510 7.680 ;
        RECT 82.960 7.600 83.260 7.680 ;
        RECT 88.710 7.600 89.010 7.680 ;
    END
  END RWL[12]
  PIN WWL[12]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 7.420 4.730 7.540 ;
        RECT 10.190 7.420 10.480 7.540 ;
        RECT 15.940 7.420 16.230 7.540 ;
        RECT 21.690 7.420 21.980 7.540 ;
        RECT 27.440 7.420 27.730 7.540 ;
        RECT 33.190 7.420 33.480 7.540 ;
        RECT 38.940 7.420 39.230 7.540 ;
        RECT 44.690 7.420 44.980 7.540 ;
        RECT 50.440 7.420 50.730 7.540 ;
        RECT 56.190 7.420 56.480 7.540 ;
        RECT 61.940 7.420 62.230 7.540 ;
        RECT 67.690 7.420 67.980 7.540 ;
        RECT 73.440 7.420 73.730 7.540 ;
        RECT 79.190 7.420 79.480 7.540 ;
        RECT 84.940 7.420 85.230 7.540 ;
        RECT 90.690 7.420 90.980 7.540 ;
        RECT -45.490 7.280 94.660 7.420 ;
        RECT 6.050 7.160 6.340 7.280 ;
        RECT 11.800 7.160 12.090 7.280 ;
        RECT 17.550 7.160 17.840 7.280 ;
        RECT 23.300 7.160 23.590 7.280 ;
        RECT 29.050 7.160 29.340 7.280 ;
        RECT 34.800 7.160 35.090 7.280 ;
        RECT 40.550 7.160 40.840 7.280 ;
        RECT 46.300 7.160 46.590 7.280 ;
        RECT 52.050 7.160 52.340 7.280 ;
        RECT 57.800 7.160 58.090 7.280 ;
        RECT 63.550 7.160 63.840 7.280 ;
        RECT 69.300 7.160 69.590 7.280 ;
        RECT 75.050 7.160 75.340 7.280 ;
        RECT 80.800 7.160 81.090 7.280 ;
        RECT 86.550 7.160 86.840 7.280 ;
        RECT 92.300 7.160 92.590 7.280 ;
    END
  END WWL[12]
  PIN RWLB[12]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 7.010 8.310 7.110 ;
        RECT 13.760 7.010 14.060 7.110 ;
        RECT 19.510 7.010 19.810 7.110 ;
        RECT 25.260 7.010 25.560 7.110 ;
        RECT 31.010 7.010 31.310 7.110 ;
        RECT 36.760 7.010 37.060 7.110 ;
        RECT 42.510 7.010 42.810 7.110 ;
        RECT 48.260 7.010 48.560 7.110 ;
        RECT 54.010 7.010 54.310 7.110 ;
        RECT 59.760 7.010 60.060 7.110 ;
        RECT 65.510 7.010 65.810 7.110 ;
        RECT 71.260 7.010 71.560 7.110 ;
        RECT 77.010 7.010 77.310 7.110 ;
        RECT 82.760 7.010 83.060 7.110 ;
        RECT 88.510 7.010 88.810 7.110 ;
        RECT 94.260 7.010 94.560 7.110 ;
        RECT -45.490 6.870 94.660 7.010 ;
        RECT 8.010 6.780 8.310 6.870 ;
        RECT 13.760 6.780 14.060 6.870 ;
        RECT 19.510 6.780 19.810 6.870 ;
        RECT 25.260 6.780 25.560 6.870 ;
        RECT 31.010 6.780 31.310 6.870 ;
        RECT 36.760 6.780 37.060 6.870 ;
        RECT 42.510 6.780 42.810 6.870 ;
        RECT 48.260 6.780 48.560 6.870 ;
        RECT 54.010 6.780 54.310 6.870 ;
        RECT 59.760 6.780 60.060 6.870 ;
        RECT 65.510 6.780 65.810 6.870 ;
        RECT 71.260 6.780 71.560 6.870 ;
        RECT 77.010 6.780 77.310 6.870 ;
        RECT 82.760 6.780 83.060 6.870 ;
        RECT 88.510 6.780 88.810 6.870 ;
        RECT 94.260 6.780 94.560 6.870 ;
    END
  END RWLB[12]
  PIN RWL[13]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 5.410 2.760 5.480 ;
        RECT 8.210 5.410 8.510 5.480 ;
        RECT 13.960 5.410 14.260 5.480 ;
        RECT 19.710 5.410 20.010 5.480 ;
        RECT 25.460 5.410 25.760 5.480 ;
        RECT 31.210 5.410 31.510 5.480 ;
        RECT 36.960 5.410 37.260 5.480 ;
        RECT 42.710 5.410 43.010 5.480 ;
        RECT 48.460 5.410 48.760 5.480 ;
        RECT 54.210 5.410 54.510 5.480 ;
        RECT 59.960 5.410 60.260 5.480 ;
        RECT 65.710 5.410 66.010 5.480 ;
        RECT 71.460 5.410 71.760 5.480 ;
        RECT 77.210 5.410 77.510 5.480 ;
        RECT 82.960 5.410 83.260 5.480 ;
        RECT 88.710 5.410 89.010 5.480 ;
        RECT -45.490 5.270 94.660 5.410 ;
        RECT 2.460 5.190 2.760 5.270 ;
        RECT 8.210 5.190 8.510 5.270 ;
        RECT 13.960 5.190 14.260 5.270 ;
        RECT 19.710 5.190 20.010 5.270 ;
        RECT 25.460 5.190 25.760 5.270 ;
        RECT 31.210 5.190 31.510 5.270 ;
        RECT 36.960 5.190 37.260 5.270 ;
        RECT 42.710 5.190 43.010 5.270 ;
        RECT 48.460 5.190 48.760 5.270 ;
        RECT 54.210 5.190 54.510 5.270 ;
        RECT 59.960 5.190 60.260 5.270 ;
        RECT 65.710 5.190 66.010 5.270 ;
        RECT 71.460 5.190 71.760 5.270 ;
        RECT 77.210 5.190 77.510 5.270 ;
        RECT 82.960 5.190 83.260 5.270 ;
        RECT 88.710 5.190 89.010 5.270 ;
    END
  END RWL[13]
  PIN WWL[13]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 5.010 4.730 5.130 ;
        RECT 10.190 5.010 10.480 5.130 ;
        RECT 15.940 5.010 16.230 5.130 ;
        RECT 21.690 5.010 21.980 5.130 ;
        RECT 27.440 5.010 27.730 5.130 ;
        RECT 33.190 5.010 33.480 5.130 ;
        RECT 38.940 5.010 39.230 5.130 ;
        RECT 44.690 5.010 44.980 5.130 ;
        RECT 50.440 5.010 50.730 5.130 ;
        RECT 56.190 5.010 56.480 5.130 ;
        RECT 61.940 5.010 62.230 5.130 ;
        RECT 67.690 5.010 67.980 5.130 ;
        RECT 73.440 5.010 73.730 5.130 ;
        RECT 79.190 5.010 79.480 5.130 ;
        RECT 84.940 5.010 85.230 5.130 ;
        RECT 90.690 5.010 90.980 5.130 ;
        RECT -45.490 4.870 94.660 5.010 ;
        RECT 6.050 4.750 6.340 4.870 ;
        RECT 11.800 4.750 12.090 4.870 ;
        RECT 17.550 4.750 17.840 4.870 ;
        RECT 23.300 4.750 23.590 4.870 ;
        RECT 29.050 4.750 29.340 4.870 ;
        RECT 34.800 4.750 35.090 4.870 ;
        RECT 40.550 4.750 40.840 4.870 ;
        RECT 46.300 4.750 46.590 4.870 ;
        RECT 52.050 4.750 52.340 4.870 ;
        RECT 57.800 4.750 58.090 4.870 ;
        RECT 63.550 4.750 63.840 4.870 ;
        RECT 69.300 4.750 69.590 4.870 ;
        RECT 75.050 4.750 75.340 4.870 ;
        RECT 80.800 4.750 81.090 4.870 ;
        RECT 86.550 4.750 86.840 4.870 ;
        RECT 92.300 4.750 92.590 4.870 ;
    END
  END WWL[13]
  PIN RWLB[13]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 4.600 8.310 4.700 ;
        RECT 13.760 4.600 14.060 4.700 ;
        RECT 19.510 4.600 19.810 4.700 ;
        RECT 25.260 4.600 25.560 4.700 ;
        RECT 31.010 4.600 31.310 4.700 ;
        RECT 36.760 4.600 37.060 4.700 ;
        RECT 42.510 4.600 42.810 4.700 ;
        RECT 48.260 4.600 48.560 4.700 ;
        RECT 54.010 4.600 54.310 4.700 ;
        RECT 59.760 4.600 60.060 4.700 ;
        RECT 65.510 4.600 65.810 4.700 ;
        RECT 71.260 4.600 71.560 4.700 ;
        RECT 77.010 4.600 77.310 4.700 ;
        RECT 82.760 4.600 83.060 4.700 ;
        RECT 88.510 4.600 88.810 4.700 ;
        RECT 94.260 4.600 94.560 4.700 ;
        RECT -45.490 4.460 94.660 4.600 ;
        RECT 8.010 4.370 8.310 4.460 ;
        RECT 13.760 4.370 14.060 4.460 ;
        RECT 19.510 4.370 19.810 4.460 ;
        RECT 25.260 4.370 25.560 4.460 ;
        RECT 31.010 4.370 31.310 4.460 ;
        RECT 36.760 4.370 37.060 4.460 ;
        RECT 42.510 4.370 42.810 4.460 ;
        RECT 48.260 4.370 48.560 4.460 ;
        RECT 54.010 4.370 54.310 4.460 ;
        RECT 59.760 4.370 60.060 4.460 ;
        RECT 65.510 4.370 65.810 4.460 ;
        RECT 71.260 4.370 71.560 4.460 ;
        RECT 77.010 4.370 77.310 4.460 ;
        RECT 82.760 4.370 83.060 4.460 ;
        RECT 88.510 4.370 88.810 4.460 ;
        RECT 94.260 4.370 94.560 4.460 ;
    END
  END RWLB[13]
  PIN RWL[14]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 3.000 2.760 3.070 ;
        RECT 8.210 3.000 8.510 3.070 ;
        RECT 13.960 3.000 14.260 3.070 ;
        RECT 19.710 3.000 20.010 3.070 ;
        RECT 25.460 3.000 25.760 3.070 ;
        RECT 31.210 3.000 31.510 3.070 ;
        RECT 36.960 3.000 37.260 3.070 ;
        RECT 42.710 3.000 43.010 3.070 ;
        RECT 48.460 3.000 48.760 3.070 ;
        RECT 54.210 3.000 54.510 3.070 ;
        RECT 59.960 3.000 60.260 3.070 ;
        RECT 65.710 3.000 66.010 3.070 ;
        RECT 71.460 3.000 71.760 3.070 ;
        RECT 77.210 3.000 77.510 3.070 ;
        RECT 82.960 3.000 83.260 3.070 ;
        RECT 88.710 3.000 89.010 3.070 ;
        RECT -45.490 2.860 94.660 3.000 ;
        RECT 2.460 2.780 2.760 2.860 ;
        RECT 8.210 2.780 8.510 2.860 ;
        RECT 13.960 2.780 14.260 2.860 ;
        RECT 19.710 2.780 20.010 2.860 ;
        RECT 25.460 2.780 25.760 2.860 ;
        RECT 31.210 2.780 31.510 2.860 ;
        RECT 36.960 2.780 37.260 2.860 ;
        RECT 42.710 2.780 43.010 2.860 ;
        RECT 48.460 2.780 48.760 2.860 ;
        RECT 54.210 2.780 54.510 2.860 ;
        RECT 59.960 2.780 60.260 2.860 ;
        RECT 65.710 2.780 66.010 2.860 ;
        RECT 71.460 2.780 71.760 2.860 ;
        RECT 77.210 2.780 77.510 2.860 ;
        RECT 82.960 2.780 83.260 2.860 ;
        RECT 88.710 2.780 89.010 2.860 ;
    END
  END RWL[14]
  PIN WWL[14]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 2.600 4.730 2.720 ;
        RECT 10.190 2.600 10.480 2.720 ;
        RECT 15.940 2.600 16.230 2.720 ;
        RECT 21.690 2.600 21.980 2.720 ;
        RECT 27.440 2.600 27.730 2.720 ;
        RECT 33.190 2.600 33.480 2.720 ;
        RECT 38.940 2.600 39.230 2.720 ;
        RECT 44.690 2.600 44.980 2.720 ;
        RECT 50.440 2.600 50.730 2.720 ;
        RECT 56.190 2.600 56.480 2.720 ;
        RECT 61.940 2.600 62.230 2.720 ;
        RECT 67.690 2.600 67.980 2.720 ;
        RECT 73.440 2.600 73.730 2.720 ;
        RECT 79.190 2.600 79.480 2.720 ;
        RECT 84.940 2.600 85.230 2.720 ;
        RECT 90.690 2.600 90.980 2.720 ;
        RECT -45.490 2.460 94.660 2.600 ;
        RECT 6.050 2.340 6.340 2.460 ;
        RECT 11.800 2.340 12.090 2.460 ;
        RECT 17.550 2.340 17.840 2.460 ;
        RECT 23.300 2.340 23.590 2.460 ;
        RECT 29.050 2.340 29.340 2.460 ;
        RECT 34.800 2.340 35.090 2.460 ;
        RECT 40.550 2.340 40.840 2.460 ;
        RECT 46.300 2.340 46.590 2.460 ;
        RECT 52.050 2.340 52.340 2.460 ;
        RECT 57.800 2.340 58.090 2.460 ;
        RECT 63.550 2.340 63.840 2.460 ;
        RECT 69.300 2.340 69.590 2.460 ;
        RECT 75.050 2.340 75.340 2.460 ;
        RECT 80.800 2.340 81.090 2.460 ;
        RECT 86.550 2.340 86.840 2.460 ;
        RECT 92.300 2.340 92.590 2.460 ;
    END
  END WWL[14]
  PIN RWLB[14]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 2.190 8.310 2.290 ;
        RECT 13.760 2.190 14.060 2.290 ;
        RECT 19.510 2.190 19.810 2.290 ;
        RECT 25.260 2.190 25.560 2.290 ;
        RECT 31.010 2.190 31.310 2.290 ;
        RECT 36.760 2.190 37.060 2.290 ;
        RECT 42.510 2.190 42.810 2.290 ;
        RECT 48.260 2.190 48.560 2.290 ;
        RECT 54.010 2.190 54.310 2.290 ;
        RECT 59.760 2.190 60.060 2.290 ;
        RECT 65.510 2.190 65.810 2.290 ;
        RECT 71.260 2.190 71.560 2.290 ;
        RECT 77.010 2.190 77.310 2.290 ;
        RECT 82.760 2.190 83.060 2.290 ;
        RECT 88.510 2.190 88.810 2.290 ;
        RECT 94.260 2.190 94.560 2.290 ;
        RECT -45.490 2.050 94.660 2.190 ;
        RECT 8.010 1.960 8.310 2.050 ;
        RECT 13.760 1.960 14.060 2.050 ;
        RECT 19.510 1.960 19.810 2.050 ;
        RECT 25.260 1.960 25.560 2.050 ;
        RECT 31.010 1.960 31.310 2.050 ;
        RECT 36.760 1.960 37.060 2.050 ;
        RECT 42.510 1.960 42.810 2.050 ;
        RECT 48.260 1.960 48.560 2.050 ;
        RECT 54.010 1.960 54.310 2.050 ;
        RECT 59.760 1.960 60.060 2.050 ;
        RECT 65.510 1.960 65.810 2.050 ;
        RECT 71.260 1.960 71.560 2.050 ;
        RECT 77.010 1.960 77.310 2.050 ;
        RECT 82.760 1.960 83.060 2.050 ;
        RECT 88.510 1.960 88.810 2.050 ;
        RECT 94.260 1.960 94.560 2.050 ;
    END
  END RWLB[14]
  PIN RWL[15]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 2.460 0.590 2.760 0.660 ;
        RECT 8.210 0.590 8.510 0.660 ;
        RECT 13.960 0.590 14.260 0.660 ;
        RECT 19.710 0.590 20.010 0.660 ;
        RECT 25.460 0.590 25.760 0.660 ;
        RECT 31.210 0.590 31.510 0.660 ;
        RECT 36.960 0.590 37.260 0.660 ;
        RECT 42.710 0.590 43.010 0.660 ;
        RECT 48.460 0.590 48.760 0.660 ;
        RECT 54.210 0.590 54.510 0.660 ;
        RECT 59.960 0.590 60.260 0.660 ;
        RECT 65.710 0.590 66.010 0.660 ;
        RECT 71.460 0.590 71.760 0.660 ;
        RECT 77.210 0.590 77.510 0.660 ;
        RECT 82.960 0.590 83.260 0.660 ;
        RECT 88.710 0.590 89.010 0.660 ;
        RECT -45.490 0.450 94.660 0.590 ;
        RECT 2.460 0.370 2.760 0.450 ;
        RECT 8.210 0.370 8.510 0.450 ;
        RECT 13.960 0.370 14.260 0.450 ;
        RECT 19.710 0.370 20.010 0.450 ;
        RECT 25.460 0.370 25.760 0.450 ;
        RECT 31.210 0.370 31.510 0.450 ;
        RECT 36.960 0.370 37.260 0.450 ;
        RECT 42.710 0.370 43.010 0.450 ;
        RECT 48.460 0.370 48.760 0.450 ;
        RECT 54.210 0.370 54.510 0.450 ;
        RECT 59.960 0.370 60.260 0.450 ;
        RECT 65.710 0.370 66.010 0.450 ;
        RECT 71.460 0.370 71.760 0.450 ;
        RECT 77.210 0.370 77.510 0.450 ;
        RECT 82.960 0.370 83.260 0.450 ;
        RECT 88.710 0.370 89.010 0.450 ;
    END
  END RWL[15]
  PIN WWL[15]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 0.190 4.730 0.310 ;
        RECT 10.190 0.190 10.480 0.310 ;
        RECT 15.940 0.190 16.230 0.310 ;
        RECT 21.690 0.190 21.980 0.310 ;
        RECT 27.440 0.190 27.730 0.310 ;
        RECT 33.190 0.190 33.480 0.310 ;
        RECT 38.940 0.190 39.230 0.310 ;
        RECT 44.690 0.190 44.980 0.310 ;
        RECT 50.440 0.190 50.730 0.310 ;
        RECT 56.190 0.190 56.480 0.310 ;
        RECT 61.940 0.190 62.230 0.310 ;
        RECT 67.690 0.190 67.980 0.310 ;
        RECT 73.440 0.190 73.730 0.310 ;
        RECT 79.190 0.190 79.480 0.310 ;
        RECT 84.940 0.190 85.230 0.310 ;
        RECT 90.690 0.190 90.980 0.310 ;
        RECT -45.490 0.050 94.660 0.190 ;
        RECT 6.050 -0.070 6.340 0.050 ;
        RECT 11.800 -0.070 12.090 0.050 ;
        RECT 17.550 -0.070 17.840 0.050 ;
        RECT 23.300 -0.070 23.590 0.050 ;
        RECT 29.050 -0.070 29.340 0.050 ;
        RECT 34.800 -0.070 35.090 0.050 ;
        RECT 40.550 -0.070 40.840 0.050 ;
        RECT 46.300 -0.070 46.590 0.050 ;
        RECT 52.050 -0.070 52.340 0.050 ;
        RECT 57.800 -0.070 58.090 0.050 ;
        RECT 63.550 -0.070 63.840 0.050 ;
        RECT 69.300 -0.070 69.590 0.050 ;
        RECT 75.050 -0.070 75.340 0.050 ;
        RECT 80.800 -0.070 81.090 0.050 ;
        RECT 86.550 -0.070 86.840 0.050 ;
        RECT 92.300 -0.070 92.590 0.050 ;
    END
  END WWL[15]
  PIN RWLB[15]
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met1 ;
        RECT 8.010 -0.220 8.310 -0.120 ;
        RECT 13.760 -0.220 14.060 -0.120 ;
        RECT 19.510 -0.220 19.810 -0.120 ;
        RECT 25.260 -0.220 25.560 -0.120 ;
        RECT 31.010 -0.220 31.310 -0.120 ;
        RECT 36.760 -0.220 37.060 -0.120 ;
        RECT 42.510 -0.220 42.810 -0.120 ;
        RECT 48.260 -0.220 48.560 -0.120 ;
        RECT 54.010 -0.220 54.310 -0.120 ;
        RECT 59.760 -0.220 60.060 -0.120 ;
        RECT 65.510 -0.220 65.810 -0.120 ;
        RECT 71.260 -0.220 71.560 -0.120 ;
        RECT 77.010 -0.220 77.310 -0.120 ;
        RECT 82.760 -0.220 83.060 -0.120 ;
        RECT 88.510 -0.220 88.810 -0.120 ;
        RECT 94.260 -0.220 94.560 -0.120 ;
        RECT -45.490 -0.360 94.660 -0.220 ;
        RECT 8.010 -0.450 8.310 -0.360 ;
        RECT 13.760 -0.450 14.060 -0.360 ;
        RECT 19.510 -0.450 19.810 -0.360 ;
        RECT 25.260 -0.450 25.560 -0.360 ;
        RECT 31.010 -0.450 31.310 -0.360 ;
        RECT 36.760 -0.450 37.060 -0.360 ;
        RECT 42.510 -0.450 42.810 -0.360 ;
        RECT 48.260 -0.450 48.560 -0.360 ;
        RECT 54.010 -0.450 54.310 -0.360 ;
        RECT 59.760 -0.450 60.060 -0.360 ;
        RECT 65.510 -0.450 65.810 -0.360 ;
        RECT 71.260 -0.450 71.560 -0.360 ;
        RECT 77.010 -0.450 77.310 -0.360 ;
        RECT 82.760 -0.450 83.060 -0.360 ;
        RECT 88.510 -0.450 88.810 -0.360 ;
        RECT 94.260 -0.450 94.560 -0.360 ;
    END
  END RWLB[15]
  PIN PRE_VLSA
    ANTENNAGATEAREA 16.799999 ;
    PORT
      LAYER met2 ;
        RECT 3.330 -14.570 3.660 -14.240 ;
        RECT 7.120 -14.570 7.440 -14.240 ;
        RECT 9.080 -14.570 9.410 -14.240 ;
        RECT 12.870 -14.570 13.190 -14.240 ;
        RECT 14.830 -14.570 15.160 -14.240 ;
        RECT 18.620 -14.570 18.940 -14.240 ;
        RECT 20.580 -14.570 20.910 -14.240 ;
        RECT 24.370 -14.570 24.690 -14.240 ;
        RECT 26.330 -14.570 26.660 -14.240 ;
        RECT 30.120 -14.570 30.440 -14.240 ;
        RECT 32.080 -14.570 32.410 -14.240 ;
        RECT 35.870 -14.570 36.190 -14.240 ;
        RECT 37.830 -14.570 38.160 -14.240 ;
        RECT 41.620 -14.570 41.940 -14.240 ;
        RECT 43.580 -14.570 43.910 -14.240 ;
        RECT 47.370 -14.570 47.690 -14.240 ;
        RECT 49.330 -14.570 49.660 -14.240 ;
        RECT 53.120 -14.570 53.440 -14.240 ;
        RECT 55.080 -14.570 55.410 -14.240 ;
        RECT 58.870 -14.570 59.190 -14.240 ;
        RECT 60.830 -14.570 61.160 -14.240 ;
        RECT 64.620 -14.570 64.940 -14.240 ;
        RECT 66.580 -14.570 66.910 -14.240 ;
        RECT 70.370 -14.570 70.690 -14.240 ;
        RECT 72.330 -14.570 72.660 -14.240 ;
        RECT 76.120 -14.570 76.440 -14.240 ;
        RECT 78.080 -14.570 78.410 -14.240 ;
        RECT 81.870 -14.570 82.190 -14.240 ;
        RECT 83.830 -14.570 84.160 -14.240 ;
        RECT 87.620 -14.570 87.940 -14.240 ;
        RECT 89.580 -14.570 89.910 -14.240 ;
        RECT 93.370 -14.570 93.690 -14.240 ;
        RECT 3.420 -18.440 3.560 -14.570 ;
        RECT 3.400 -18.770 3.730 -18.440 ;
        RECT 7.220 -18.450 7.360 -14.570 ;
        RECT 9.170 -18.440 9.310 -14.570 ;
        RECT 7.080 -18.780 7.410 -18.450 ;
        RECT 9.150 -18.770 9.480 -18.440 ;
        RECT 12.970 -18.450 13.110 -14.570 ;
        RECT 14.920 -18.440 15.060 -14.570 ;
        RECT 12.830 -18.780 13.160 -18.450 ;
        RECT 14.900 -18.770 15.230 -18.440 ;
        RECT 18.720 -18.450 18.860 -14.570 ;
        RECT 20.670 -18.440 20.810 -14.570 ;
        RECT 18.580 -18.780 18.910 -18.450 ;
        RECT 20.650 -18.770 20.980 -18.440 ;
        RECT 24.470 -18.450 24.610 -14.570 ;
        RECT 26.420 -18.440 26.560 -14.570 ;
        RECT 24.330 -18.780 24.660 -18.450 ;
        RECT 26.400 -18.770 26.730 -18.440 ;
        RECT 30.220 -18.450 30.360 -14.570 ;
        RECT 32.170 -18.440 32.310 -14.570 ;
        RECT 30.080 -18.780 30.410 -18.450 ;
        RECT 32.150 -18.770 32.480 -18.440 ;
        RECT 35.970 -18.450 36.110 -14.570 ;
        RECT 37.920 -18.440 38.060 -14.570 ;
        RECT 35.830 -18.780 36.160 -18.450 ;
        RECT 37.900 -18.770 38.230 -18.440 ;
        RECT 41.720 -18.450 41.860 -14.570 ;
        RECT 43.670 -18.440 43.810 -14.570 ;
        RECT 41.580 -18.780 41.910 -18.450 ;
        RECT 43.650 -18.770 43.980 -18.440 ;
        RECT 47.470 -18.450 47.610 -14.570 ;
        RECT 49.420 -18.440 49.560 -14.570 ;
        RECT 47.330 -18.780 47.660 -18.450 ;
        RECT 49.400 -18.770 49.730 -18.440 ;
        RECT 53.220 -18.450 53.360 -14.570 ;
        RECT 55.170 -18.440 55.310 -14.570 ;
        RECT 53.080 -18.780 53.410 -18.450 ;
        RECT 55.150 -18.770 55.480 -18.440 ;
        RECT 58.970 -18.450 59.110 -14.570 ;
        RECT 60.920 -18.440 61.060 -14.570 ;
        RECT 58.830 -18.780 59.160 -18.450 ;
        RECT 60.900 -18.770 61.230 -18.440 ;
        RECT 64.720 -18.450 64.860 -14.570 ;
        RECT 66.670 -18.440 66.810 -14.570 ;
        RECT 64.580 -18.780 64.910 -18.450 ;
        RECT 66.650 -18.770 66.980 -18.440 ;
        RECT 70.470 -18.450 70.610 -14.570 ;
        RECT 72.420 -18.440 72.560 -14.570 ;
        RECT 70.330 -18.780 70.660 -18.450 ;
        RECT 72.400 -18.770 72.730 -18.440 ;
        RECT 76.220 -18.450 76.360 -14.570 ;
        RECT 78.170 -18.440 78.310 -14.570 ;
        RECT 76.080 -18.780 76.410 -18.450 ;
        RECT 78.150 -18.770 78.480 -18.440 ;
        RECT 81.970 -18.450 82.110 -14.570 ;
        RECT 83.920 -18.440 84.060 -14.570 ;
        RECT 81.830 -18.780 82.160 -18.450 ;
        RECT 83.900 -18.770 84.230 -18.440 ;
        RECT 87.720 -18.450 87.860 -14.570 ;
        RECT 89.670 -18.440 89.810 -14.570 ;
        RECT 87.580 -18.780 87.910 -18.450 ;
        RECT 89.650 -18.770 89.980 -18.440 ;
        RECT 93.470 -18.450 93.610 -14.570 ;
        RECT 93.330 -18.780 93.660 -18.450 ;
    END
  END PRE_VLSA
  PIN WE
    ANTENNAGATEAREA 4.800000 ;
    PORT
      LAYER met1 ;
        RECT 4.270 -19.500 4.600 -19.440 ;
        RECT 6.150 -19.500 6.480 -19.440 ;
        RECT 10.020 -19.500 10.350 -19.440 ;
        RECT 11.900 -19.500 12.230 -19.440 ;
        RECT 15.770 -19.500 16.100 -19.440 ;
        RECT 17.650 -19.500 17.980 -19.440 ;
        RECT 21.520 -19.500 21.850 -19.440 ;
        RECT 23.400 -19.500 23.730 -19.440 ;
        RECT 27.270 -19.500 27.600 -19.440 ;
        RECT 29.150 -19.500 29.480 -19.440 ;
        RECT 33.020 -19.500 33.350 -19.440 ;
        RECT 34.900 -19.500 35.230 -19.440 ;
        RECT 38.770 -19.500 39.100 -19.440 ;
        RECT 40.650 -19.500 40.980 -19.440 ;
        RECT 44.520 -19.500 44.850 -19.440 ;
        RECT 46.400 -19.500 46.730 -19.440 ;
        RECT 50.270 -19.500 50.600 -19.440 ;
        RECT 52.150 -19.500 52.480 -19.440 ;
        RECT 56.020 -19.500 56.350 -19.440 ;
        RECT 57.900 -19.500 58.230 -19.440 ;
        RECT 61.770 -19.500 62.100 -19.440 ;
        RECT 63.650 -19.500 63.980 -19.440 ;
        RECT 67.520 -19.500 67.850 -19.440 ;
        RECT 69.400 -19.500 69.730 -19.440 ;
        RECT 73.270 -19.500 73.600 -19.440 ;
        RECT 75.150 -19.500 75.480 -19.440 ;
        RECT 79.020 -19.500 79.350 -19.440 ;
        RECT 80.900 -19.500 81.230 -19.440 ;
        RECT 84.770 -19.500 85.100 -19.440 ;
        RECT 86.650 -19.500 86.980 -19.440 ;
        RECT 90.520 -19.500 90.850 -19.440 ;
        RECT 92.400 -19.500 92.730 -19.440 ;
        RECT -45.490 -19.640 94.660 -19.500 ;
        RECT 4.270 -19.690 4.600 -19.640 ;
        RECT 6.150 -19.690 6.480 -19.640 ;
        RECT 10.020 -19.690 10.350 -19.640 ;
        RECT 11.900 -19.690 12.230 -19.640 ;
        RECT 15.770 -19.690 16.100 -19.640 ;
        RECT 17.650 -19.690 17.980 -19.640 ;
        RECT 21.520 -19.690 21.850 -19.640 ;
        RECT 23.400 -19.690 23.730 -19.640 ;
        RECT 27.270 -19.690 27.600 -19.640 ;
        RECT 29.150 -19.690 29.480 -19.640 ;
        RECT 33.020 -19.690 33.350 -19.640 ;
        RECT 34.900 -19.690 35.230 -19.640 ;
        RECT 38.770 -19.690 39.100 -19.640 ;
        RECT 40.650 -19.690 40.980 -19.640 ;
        RECT 44.520 -19.690 44.850 -19.640 ;
        RECT 46.400 -19.690 46.730 -19.640 ;
        RECT 50.270 -19.690 50.600 -19.640 ;
        RECT 52.150 -19.690 52.480 -19.640 ;
        RECT 56.020 -19.690 56.350 -19.640 ;
        RECT 57.900 -19.690 58.230 -19.640 ;
        RECT 61.770 -19.690 62.100 -19.640 ;
        RECT 63.650 -19.690 63.980 -19.640 ;
        RECT 67.520 -19.690 67.850 -19.640 ;
        RECT 69.400 -19.690 69.730 -19.640 ;
        RECT 73.270 -19.690 73.600 -19.640 ;
        RECT 75.150 -19.690 75.480 -19.640 ;
        RECT 79.020 -19.690 79.350 -19.640 ;
        RECT 80.900 -19.690 81.230 -19.640 ;
        RECT 84.770 -19.690 85.100 -19.640 ;
        RECT 86.650 -19.690 86.980 -19.640 ;
        RECT 90.520 -19.690 90.850 -19.640 ;
        RECT 92.400 -19.690 92.730 -19.640 ;
    END
  END WE
  PIN PRE_CLSA
    ANTENNAGATEAREA 76.799995 ;
    PORT
      LAYER met2 ;
        RECT -39.880 -31.540 -39.620 -31.220 ;
        RECT -39.820 -58.540 -39.680 -31.540 ;
        RECT -39.870 -58.860 -39.610 -58.540 ;
        RECT -39.820 -85.870 -39.680 -58.860 ;
        RECT -39.910 -86.190 -39.590 -85.870 ;
        RECT -39.820 -90.250 -39.680 -86.190 ;
    END
  END PRE_CLSA
  PIN VCLP
    ANTENNAGATEAREA 134.399994 ;
    PORT
      LAYER met2 ;
        RECT -40.540 -36.570 -40.280 -36.250 ;
        RECT -40.480 -53.510 -40.340 -36.570 ;
        RECT -40.540 -53.830 -40.280 -53.510 ;
        RECT -40.480 -63.580 -40.340 -53.830 ;
        RECT -40.570 -63.900 -40.250 -63.580 ;
        RECT -40.480 -80.840 -40.340 -63.900 ;
        RECT -40.570 -81.160 -40.250 -80.840 ;
        RECT -40.480 -90.250 -40.340 -81.160 ;
    END
  END VCLP
  PIN SAEN
    ANTENNAGATEAREA 9.240000 ;
    PORT
      LAYER met2 ;
        RECT -41.200 -36.970 -40.940 -36.650 ;
        RECT -41.140 -53.110 -41.000 -36.970 ;
        RECT -41.230 -53.430 -40.910 -53.110 ;
        RECT -41.140 -63.980 -41.000 -53.430 ;
        RECT -41.230 -64.300 -40.910 -63.980 ;
        RECT -41.140 -80.440 -41.000 -64.300 ;
        RECT -41.230 -80.760 -40.910 -80.440 ;
        RECT -41.140 -90.250 -41.000 -80.760 ;
    END
  END SAEN
  PIN ADC0_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -31.480 -36.130 -31.220 -35.810 ;
        RECT -31.420 -90.170 -31.280 -36.130 ;
    END
  END ADC0_OUT[0]
  PIN ADC0_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -31.070 -54.260 -30.810 -53.940 ;
        RECT -31.010 -90.170 -30.870 -54.260 ;
    END
  END ADC0_OUT[1]
  PIN ADC0_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -30.670 -63.460 -30.410 -63.140 ;
        RECT -30.610 -90.170 -30.470 -63.460 ;
    END
  END ADC0_OUT[2]
  PIN ADC0_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -30.260 -81.590 -30.000 -81.270 ;
        RECT -30.200 -90.170 -30.060 -81.590 ;
    END
  END ADC0_OUT[3]
  PIN ADC1_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -19.930 -36.130 -19.670 -35.810 ;
        RECT -19.870 -90.090 -19.730 -36.130 ;
    END
  END ADC1_OUT[0]
  PIN ADC1_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -19.530 -54.260 -19.270 -53.940 ;
        RECT -19.470 -90.090 -19.330 -54.260 ;
    END
  END ADC1_OUT[1]
  PIN ADC1_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -19.140 -63.460 -18.820 -63.140 ;
        RECT -19.050 -90.090 -18.910 -63.460 ;
    END
  END ADC1_OUT[2]
  PIN ADC1_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -18.700 -81.590 -18.440 -81.270 ;
        RECT -18.640 -90.090 -18.500 -81.590 ;
    END
  END ADC1_OUT[3]
  PIN ADC2_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -8.240 -36.130 -7.980 -35.810 ;
        RECT -8.180 -89.860 -8.040 -36.130 ;
    END
  END ADC2_OUT[0]
  PIN ADC2_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -7.840 -54.260 -7.580 -53.940 ;
        RECT -7.780 -89.860 -7.640 -54.260 ;
    END
  END ADC2_OUT[1]
  PIN ADC2_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -7.450 -63.460 -7.130 -63.140 ;
        RECT -7.360 -89.860 -7.220 -63.460 ;
    END
  END ADC2_OUT[2]
  PIN ADC2_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT -7.010 -81.590 -6.750 -81.270 ;
        RECT -6.950 -89.860 -6.810 -81.590 ;
    END
  END ADC2_OUT[3]
  PIN ADC3_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 3.670 -36.130 3.930 -35.810 ;
        RECT 3.730 -89.780 3.870 -36.130 ;
    END
  END ADC3_OUT[0]
  PIN ADC3_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 4.070 -54.260 4.330 -53.940 ;
        RECT 4.130 -89.780 4.270 -54.260 ;
    END
  END ADC3_OUT[1]
  PIN ADC3_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 4.460 -63.460 4.780 -63.140 ;
        RECT 4.550 -89.780 4.690 -63.460 ;
    END
  END ADC3_OUT[2]
  PIN ADC3_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 4.900 -81.590 5.160 -81.270 ;
        RECT 4.960 -89.780 5.100 -81.590 ;
    END
  END ADC3_OUT[3]
  PIN ADC4_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 15.440 -36.130 15.700 -35.810 ;
        RECT 15.500 -89.950 15.640 -36.130 ;
    END
  END ADC4_OUT[0]
  PIN ADC4_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 15.840 -54.260 16.100 -53.940 ;
        RECT 15.900 -89.950 16.040 -54.260 ;
    END
  END ADC4_OUT[1]
  PIN ADC4_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 16.230 -63.460 16.550 -63.140 ;
        RECT 16.320 -89.950 16.460 -63.460 ;
    END
  END ADC4_OUT[2]
  PIN ADC4_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 16.670 -81.590 16.930 -81.270 ;
        RECT 16.730 -89.950 16.870 -81.590 ;
    END
  END ADC4_OUT[3]
  PIN ADC5_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 27.210 -36.130 27.470 -35.810 ;
        RECT 27.270 -90.070 27.410 -36.130 ;
    END
  END ADC5_OUT[0]
  PIN ADC5_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 27.610 -54.260 27.870 -53.940 ;
        RECT 27.670 -90.070 27.810 -54.260 ;
    END
  END ADC5_OUT[1]
  PIN ADC5_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 28.000 -63.460 28.320 -63.140 ;
        RECT 28.090 -90.070 28.230 -63.460 ;
    END
  END ADC5_OUT[2]
  PIN ADC5_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 28.440 -81.590 28.700 -81.270 ;
        RECT 28.500 -90.070 28.640 -81.590 ;
    END
  END ADC5_OUT[3]
  PIN ADC6_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 39.030 -36.130 39.290 -35.810 ;
        RECT 39.090 -90.180 39.230 -36.130 ;
    END
  END ADC6_OUT[0]
  PIN ADC6_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 39.430 -54.260 39.690 -53.940 ;
        RECT 39.490 -90.180 39.630 -54.260 ;
    END
  END ADC6_OUT[1]
  PIN ADC6_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 39.820 -63.460 40.140 -63.140 ;
        RECT 39.910 -90.180 40.050 -63.460 ;
    END
  END ADC6_OUT[2]
  PIN ADC6_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 40.260 -81.590 40.520 -81.270 ;
        RECT 40.320 -90.180 40.460 -81.590 ;
    END
  END ADC6_OUT[3]
  PIN ADC7_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 50.890 -36.130 51.150 -35.810 ;
        RECT 50.950 -90.260 51.090 -36.130 ;
    END
  END ADC7_OUT[0]
  PIN ADC7_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 51.290 -54.260 51.550 -53.940 ;
        RECT 51.350 -90.260 51.490 -54.260 ;
    END
  END ADC7_OUT[1]
  PIN ADC7_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 51.680 -63.460 52.000 -63.140 ;
        RECT 51.770 -90.260 51.910 -63.460 ;
    END
  END ADC7_OUT[2]
  PIN ADC7_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 52.120 -81.590 52.380 -81.270 ;
        RECT 52.180 -90.260 52.320 -81.590 ;
    END
  END ADC7_OUT[3]
  PIN ADC8_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 62.680 -36.130 62.940 -35.810 ;
        RECT 62.740 -90.230 62.880 -36.130 ;
    END
  END ADC8_OUT[0]
  PIN ADC8_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 63.080 -54.260 63.340 -53.940 ;
        RECT 63.140 -90.230 63.280 -54.260 ;
    END
  END ADC8_OUT[1]
  PIN ADC8_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 63.470 -63.460 63.790 -63.140 ;
        RECT 63.560 -90.230 63.700 -63.460 ;
    END
  END ADC8_OUT[2]
  PIN ADC8_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 63.910 -81.590 64.170 -81.270 ;
        RECT 63.970 -90.230 64.110 -81.590 ;
    END
  END ADC8_OUT[3]
  PIN ADC9_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 74.560 -36.130 74.820 -35.810 ;
        RECT 74.620 -90.120 74.760 -36.130 ;
    END
  END ADC9_OUT[0]
  PIN ADC9_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 74.960 -54.260 75.220 -53.940 ;
        RECT 75.020 -90.120 75.160 -54.260 ;
    END
  END ADC9_OUT[1]
  PIN ADC9_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 75.350 -63.460 75.670 -63.140 ;
        RECT 75.440 -90.120 75.580 -63.460 ;
    END
  END ADC9_OUT[2]
  PIN ADC9_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 75.790 -81.590 76.050 -81.270 ;
        RECT 75.850 -90.120 75.990 -81.590 ;
    END
  END ADC9_OUT[3]
  PIN ADC10_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 86.290 -36.130 86.550 -35.810 ;
        RECT 86.350 -90.270 86.490 -36.130 ;
    END
  END ADC10_OUT[0]
  PIN ADC10_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 86.690 -54.260 86.950 -53.940 ;
        RECT 86.750 -90.270 86.890 -54.260 ;
    END
  END ADC10_OUT[1]
  PIN ADC10_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 87.080 -63.460 87.400 -63.140 ;
        RECT 87.170 -90.270 87.310 -63.460 ;
    END
  END ADC10_OUT[2]
  PIN ADC10_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 87.520 -81.590 87.780 -81.270 ;
        RECT 87.580 -90.270 87.720 -81.590 ;
    END
  END ADC10_OUT[3]
  PIN ADC11_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 98.110 -36.130 98.370 -35.810 ;
        RECT 98.170 -90.350 98.310 -36.130 ;
    END
  END ADC11_OUT[0]
  PIN ADC11_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 98.510 -54.260 98.770 -53.940 ;
        RECT 98.570 -90.350 98.710 -54.260 ;
    END
  END ADC11_OUT[1]
  PIN ADC11_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 98.900 -63.460 99.220 -63.140 ;
        RECT 98.990 -90.350 99.130 -63.460 ;
    END
  END ADC11_OUT[2]
  PIN ADC11_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 99.340 -81.590 99.600 -81.270 ;
        RECT 99.400 -90.350 99.540 -81.590 ;
    END
  END ADC11_OUT[3]
  PIN ADC12_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 110.000 -36.130 110.260 -35.810 ;
        RECT 110.060 -90.170 110.200 -36.130 ;
    END
  END ADC12_OUT[0]
  PIN ADC12_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 110.400 -54.260 110.660 -53.940 ;
        RECT 110.460 -90.170 110.600 -54.260 ;
    END
  END ADC12_OUT[1]
  PIN ADC12_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 110.790 -63.460 111.110 -63.140 ;
        RECT 110.880 -90.170 111.020 -63.460 ;
    END
  END ADC12_OUT[2]
  PIN ADC12_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 111.230 -81.590 111.490 -81.270 ;
        RECT 111.290 -90.170 111.430 -81.590 ;
    END
  END ADC12_OUT[3]
  PIN ADC13_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 121.950 -36.130 122.210 -35.810 ;
        RECT 122.010 -90.130 122.150 -36.130 ;
    END
  END ADC13_OUT[0]
  PIN ADC13_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 122.350 -54.260 122.610 -53.940 ;
        RECT 122.410 -90.130 122.550 -54.260 ;
    END
  END ADC13_OUT[1]
  PIN ADC13_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 122.740 -63.460 123.060 -63.140 ;
        RECT 122.830 -90.130 122.970 -63.460 ;
    END
  END ADC13_OUT[2]
  PIN ADC13_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 123.180 -81.590 123.440 -81.270 ;
        RECT 123.240 -90.130 123.380 -81.590 ;
    END
  END ADC13_OUT[3]
  PIN ADC14_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 133.710 -36.130 133.970 -35.810 ;
        RECT 133.770 -90.070 133.910 -36.130 ;
    END
  END ADC14_OUT[0]
  PIN ADC14_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 134.110 -54.260 134.370 -53.940 ;
        RECT 134.170 -90.070 134.310 -54.260 ;
    END
  END ADC14_OUT[1]
  PIN ADC14_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 134.500 -63.460 134.820 -63.140 ;
        RECT 134.590 -90.070 134.730 -63.460 ;
    END
  END ADC14_OUT[2]
  PIN ADC14_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 134.940 -81.590 135.200 -81.270 ;
        RECT 135.000 -90.070 135.140 -81.590 ;
    END
  END ADC14_OUT[3]
  PIN ADC15_OUT[0]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 142.750 -36.130 143.010 -35.810 ;
        RECT 142.810 -90.110 142.950 -36.130 ;
    END
  END ADC15_OUT[0]
  PIN ADC15_OUT[1]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 143.150 -54.260 143.410 -53.940 ;
        RECT 143.210 -90.110 143.350 -54.260 ;
    END
  END ADC15_OUT[1]
  PIN ADC15_OUT[2]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 143.540 -63.460 143.860 -63.140 ;
        RECT 143.630 -90.110 143.770 -63.460 ;
    END
  END ADC15_OUT[2]
  PIN ADC15_OUT[3]
    ANTENNAGATEAREA 1.800000 ;
    ANTENNADIFFAREA 4.320000 ;
    PORT
      LAYER met2 ;
        RECT 143.980 -81.590 144.240 -81.270 ;
        RECT 144.040 -90.110 144.180 -81.590 ;
    END
  END ADC15_OUT[3]
  PIN Din[0]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 2.340 -20.980 2.480 53.560 ;
        RECT 2.250 -21.300 2.570 -20.980 ;
    END
  END Din[0]
  PIN Din[1]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 8.150 -20.960 8.290 53.450 ;
        RECT 8.060 -21.280 8.380 -20.960 ;
    END
  END Din[1]
  PIN Din[2]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 13.860 -20.970 14.000 53.410 ;
        RECT 13.780 -21.290 14.100 -20.970 ;
    END
  END Din[2]
  PIN Din[3]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 19.640 -20.990 19.780 53.420 ;
        RECT 19.560 -21.310 19.880 -20.990 ;
    END
  END Din[3]
  PIN Din[4]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 25.370 -20.990 25.510 53.420 ;
        RECT 25.310 -21.310 25.630 -20.990 ;
    END
  END Din[4]
  PIN Din[5]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 31.100 -21.010 31.240 53.400 ;
        RECT 31.020 -21.330 31.340 -21.010 ;
    END
  END Din[5]
  PIN Din[6]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 36.860 -21.000 37.000 53.410 ;
        RECT 36.790 -21.320 37.110 -21.000 ;
    END
  END Din[6]
  PIN Din[7]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 42.640 -20.990 42.780 53.420 ;
        RECT 42.590 -21.310 42.910 -20.990 ;
    END
  END Din[7]
  PIN Din[8]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 48.370 -20.980 48.510 53.420 ;
        RECT 48.290 -21.300 48.610 -20.980 ;
    END
  END Din[8]
  PIN Din[9]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 54.120 -21.000 54.260 53.400 ;
        RECT 54.060 -21.320 54.380 -21.000 ;
    END
  END Din[9]
  PIN Din[10]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 59.880 -20.980 60.020 53.410 ;
        RECT 59.800 -21.300 60.120 -20.980 ;
    END
  END Din[10]
  PIN Din[11]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 65.610 -20.990 65.750 53.410 ;
        RECT 65.530 -21.310 65.850 -20.990 ;
    END
  END Din[11]
  PIN Din[12]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 71.360 -21.000 71.500 53.410 ;
        RECT 71.300 -21.320 71.620 -21.000 ;
    END
  END Din[12]
  PIN Din[13]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 77.110 -21.000 77.250 53.420 ;
        RECT 77.060 -21.320 77.380 -21.000 ;
    END
  END Din[13]
  PIN Din[14]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 82.880 -21.020 83.020 53.420 ;
        RECT 82.790 -21.340 83.110 -21.020 ;
    END
  END Din[14]
  PIN Din[15]
    ANTENNAGATEAREA 0.189000 ;
    PORT
      LAYER met2 ;
        RECT 88.630 -21.020 88.770 53.420 ;
        RECT 88.540 -21.340 88.860 -21.020 ;
    END
  END Din[15]
  PIN WWLD[0]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 47.350 4.730 47.470 ;
        RECT 10.190 47.350 10.480 47.470 ;
        RECT 15.940 47.350 16.230 47.470 ;
        RECT 21.690 47.350 21.980 47.470 ;
        RECT 27.440 47.350 27.730 47.470 ;
        RECT 33.190 47.350 33.480 47.470 ;
        RECT 38.940 47.350 39.230 47.470 ;
        RECT 44.690 47.350 44.980 47.470 ;
        RECT 50.440 47.350 50.730 47.470 ;
        RECT 56.190 47.350 56.480 47.470 ;
        RECT 61.940 47.350 62.230 47.470 ;
        RECT 67.690 47.350 67.980 47.470 ;
        RECT 73.440 47.350 73.730 47.470 ;
        RECT 79.190 47.350 79.480 47.470 ;
        RECT 84.940 47.350 85.230 47.470 ;
        RECT 90.690 47.350 90.980 47.470 ;
        RECT -45.490 47.210 94.660 47.350 ;
        RECT 6.050 47.090 6.340 47.210 ;
        RECT 11.800 47.090 12.090 47.210 ;
        RECT 17.550 47.090 17.840 47.210 ;
        RECT 23.300 47.090 23.590 47.210 ;
        RECT 29.050 47.090 29.340 47.210 ;
        RECT 34.800 47.090 35.090 47.210 ;
        RECT 40.550 47.090 40.840 47.210 ;
        RECT 46.300 47.090 46.590 47.210 ;
        RECT 52.050 47.090 52.340 47.210 ;
        RECT 57.800 47.090 58.090 47.210 ;
        RECT 63.550 47.090 63.840 47.210 ;
        RECT 69.300 47.090 69.590 47.210 ;
        RECT 75.050 47.090 75.340 47.210 ;
        RECT 80.800 47.090 81.090 47.210 ;
        RECT 86.550 47.090 86.840 47.210 ;
        RECT 92.300 47.090 92.590 47.210 ;
    END
  END WWLD[0]
  PIN WWLD[1]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 44.940 4.730 45.060 ;
        RECT 10.190 44.940 10.480 45.060 ;
        RECT 15.940 44.940 16.230 45.060 ;
        RECT 21.690 44.940 21.980 45.060 ;
        RECT 27.440 44.940 27.730 45.060 ;
        RECT 33.190 44.940 33.480 45.060 ;
        RECT 38.940 44.940 39.230 45.060 ;
        RECT 44.690 44.940 44.980 45.060 ;
        RECT 50.440 44.940 50.730 45.060 ;
        RECT 56.190 44.940 56.480 45.060 ;
        RECT 61.940 44.940 62.230 45.060 ;
        RECT 67.690 44.940 67.980 45.060 ;
        RECT 73.440 44.940 73.730 45.060 ;
        RECT 79.190 44.940 79.480 45.060 ;
        RECT 84.940 44.940 85.230 45.060 ;
        RECT 90.690 44.940 90.980 45.060 ;
        RECT -45.490 44.800 94.660 44.940 ;
        RECT 6.050 44.680 6.340 44.800 ;
        RECT 11.800 44.680 12.090 44.800 ;
        RECT 17.550 44.680 17.840 44.800 ;
        RECT 23.300 44.680 23.590 44.800 ;
        RECT 29.050 44.680 29.340 44.800 ;
        RECT 34.800 44.680 35.090 44.800 ;
        RECT 40.550 44.680 40.840 44.800 ;
        RECT 46.300 44.680 46.590 44.800 ;
        RECT 52.050 44.680 52.340 44.800 ;
        RECT 57.800 44.680 58.090 44.800 ;
        RECT 63.550 44.680 63.840 44.800 ;
        RECT 69.300 44.680 69.590 44.800 ;
        RECT 75.050 44.680 75.340 44.800 ;
        RECT 80.800 44.680 81.090 44.800 ;
        RECT 86.550 44.680 86.840 44.800 ;
        RECT 92.300 44.680 92.590 44.800 ;
    END
  END WWLD[1]
  PIN WWLD[2]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 41.970 4.730 42.090 ;
        RECT 10.190 41.970 10.480 42.090 ;
        RECT 15.940 41.970 16.230 42.090 ;
        RECT 21.690 41.970 21.980 42.090 ;
        RECT 27.440 41.970 27.730 42.090 ;
        RECT 33.190 41.970 33.480 42.090 ;
        RECT 38.940 41.970 39.230 42.090 ;
        RECT 44.690 41.970 44.980 42.090 ;
        RECT 50.440 41.970 50.730 42.090 ;
        RECT 56.190 41.970 56.480 42.090 ;
        RECT 61.940 41.970 62.230 42.090 ;
        RECT 67.690 41.970 67.980 42.090 ;
        RECT 73.440 41.970 73.730 42.090 ;
        RECT 79.190 41.970 79.480 42.090 ;
        RECT 84.940 41.970 85.230 42.090 ;
        RECT 90.690 41.970 90.980 42.090 ;
        RECT -45.490 41.830 94.660 41.970 ;
        RECT 6.050 41.710 6.340 41.830 ;
        RECT 11.800 41.710 12.090 41.830 ;
        RECT 17.550 41.710 17.840 41.830 ;
        RECT 23.300 41.710 23.590 41.830 ;
        RECT 29.050 41.710 29.340 41.830 ;
        RECT 34.800 41.710 35.090 41.830 ;
        RECT 40.550 41.710 40.840 41.830 ;
        RECT 46.300 41.710 46.590 41.830 ;
        RECT 52.050 41.710 52.340 41.830 ;
        RECT 57.800 41.710 58.090 41.830 ;
        RECT 63.550 41.710 63.840 41.830 ;
        RECT 69.300 41.710 69.590 41.830 ;
        RECT 75.050 41.710 75.340 41.830 ;
        RECT 80.800 41.710 81.090 41.830 ;
        RECT 86.550 41.710 86.840 41.830 ;
        RECT 92.300 41.710 92.590 41.830 ;
    END
  END WWLD[2]
  PIN WWLD[3]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 39.560 4.730 39.680 ;
        RECT 10.190 39.560 10.480 39.680 ;
        RECT 15.940 39.560 16.230 39.680 ;
        RECT 21.690 39.560 21.980 39.680 ;
        RECT 27.440 39.560 27.730 39.680 ;
        RECT 33.190 39.560 33.480 39.680 ;
        RECT 38.940 39.560 39.230 39.680 ;
        RECT 44.690 39.560 44.980 39.680 ;
        RECT 50.440 39.560 50.730 39.680 ;
        RECT 56.190 39.560 56.480 39.680 ;
        RECT 61.940 39.560 62.230 39.680 ;
        RECT 67.690 39.560 67.980 39.680 ;
        RECT 73.440 39.560 73.730 39.680 ;
        RECT 79.190 39.560 79.480 39.680 ;
        RECT 84.940 39.560 85.230 39.680 ;
        RECT 90.690 39.560 90.980 39.680 ;
        RECT -45.490 39.420 94.660 39.560 ;
        RECT 6.050 39.300 6.340 39.420 ;
        RECT 11.800 39.300 12.090 39.420 ;
        RECT 17.550 39.300 17.840 39.420 ;
        RECT 23.300 39.300 23.590 39.420 ;
        RECT 29.050 39.300 29.340 39.420 ;
        RECT 34.800 39.300 35.090 39.420 ;
        RECT 40.550 39.300 40.840 39.420 ;
        RECT 46.300 39.300 46.590 39.420 ;
        RECT 52.050 39.300 52.340 39.420 ;
        RECT 57.800 39.300 58.090 39.420 ;
        RECT 63.550 39.300 63.840 39.420 ;
        RECT 69.300 39.300 69.590 39.420 ;
        RECT 75.050 39.300 75.340 39.420 ;
        RECT 80.800 39.300 81.090 39.420 ;
        RECT 86.550 39.300 86.840 39.420 ;
        RECT 92.300 39.300 92.590 39.420 ;
    END
  END WWLD[3]
  PIN WWLD[4]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 -2.220 4.730 -2.100 ;
        RECT 10.190 -2.220 10.480 -2.100 ;
        RECT 15.940 -2.220 16.230 -2.100 ;
        RECT 21.690 -2.220 21.980 -2.100 ;
        RECT 27.440 -2.220 27.730 -2.100 ;
        RECT 33.190 -2.220 33.480 -2.100 ;
        RECT 38.940 -2.220 39.230 -2.100 ;
        RECT 44.690 -2.220 44.980 -2.100 ;
        RECT 50.440 -2.220 50.730 -2.100 ;
        RECT 56.190 -2.220 56.480 -2.100 ;
        RECT 61.940 -2.220 62.230 -2.100 ;
        RECT 67.690 -2.220 67.980 -2.100 ;
        RECT 73.440 -2.220 73.730 -2.100 ;
        RECT 79.190 -2.220 79.480 -2.100 ;
        RECT 84.940 -2.220 85.230 -2.100 ;
        RECT 90.690 -2.220 90.980 -2.100 ;
        RECT -45.490 -2.360 94.660 -2.220 ;
        RECT 6.050 -2.480 6.340 -2.360 ;
        RECT 11.800 -2.480 12.090 -2.360 ;
        RECT 17.550 -2.480 17.840 -2.360 ;
        RECT 23.300 -2.480 23.590 -2.360 ;
        RECT 29.050 -2.480 29.340 -2.360 ;
        RECT 34.800 -2.480 35.090 -2.360 ;
        RECT 40.550 -2.480 40.840 -2.360 ;
        RECT 46.300 -2.480 46.590 -2.360 ;
        RECT 52.050 -2.480 52.340 -2.360 ;
        RECT 57.800 -2.480 58.090 -2.360 ;
        RECT 63.550 -2.480 63.840 -2.360 ;
        RECT 69.300 -2.480 69.590 -2.360 ;
        RECT 75.050 -2.480 75.340 -2.360 ;
        RECT 80.800 -2.480 81.090 -2.360 ;
        RECT 86.550 -2.480 86.840 -2.360 ;
        RECT 92.300 -2.480 92.590 -2.360 ;
    END
  END WWLD[4]
  PIN WWLD[5]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 -4.630 4.730 -4.510 ;
        RECT 10.190 -4.630 10.480 -4.510 ;
        RECT 15.940 -4.630 16.230 -4.510 ;
        RECT 21.690 -4.630 21.980 -4.510 ;
        RECT 27.440 -4.630 27.730 -4.510 ;
        RECT 33.190 -4.630 33.480 -4.510 ;
        RECT 38.940 -4.630 39.230 -4.510 ;
        RECT 44.690 -4.630 44.980 -4.510 ;
        RECT 50.440 -4.630 50.730 -4.510 ;
        RECT 56.190 -4.630 56.480 -4.510 ;
        RECT 61.940 -4.630 62.230 -4.510 ;
        RECT 67.690 -4.630 67.980 -4.510 ;
        RECT 73.440 -4.630 73.730 -4.510 ;
        RECT 79.190 -4.630 79.480 -4.510 ;
        RECT 84.940 -4.630 85.230 -4.510 ;
        RECT 90.690 -4.630 90.980 -4.510 ;
        RECT -45.490 -4.770 94.660 -4.630 ;
        RECT 6.050 -4.890 6.340 -4.770 ;
        RECT 11.800 -4.890 12.090 -4.770 ;
        RECT 17.550 -4.890 17.840 -4.770 ;
        RECT 23.300 -4.890 23.590 -4.770 ;
        RECT 29.050 -4.890 29.340 -4.770 ;
        RECT 34.800 -4.890 35.090 -4.770 ;
        RECT 40.550 -4.890 40.840 -4.770 ;
        RECT 46.300 -4.890 46.590 -4.770 ;
        RECT 52.050 -4.890 52.340 -4.770 ;
        RECT 57.800 -4.890 58.090 -4.770 ;
        RECT 63.550 -4.890 63.840 -4.770 ;
        RECT 69.300 -4.890 69.590 -4.770 ;
        RECT 75.050 -4.890 75.340 -4.770 ;
        RECT 80.800 -4.890 81.090 -4.770 ;
        RECT 86.550 -4.890 86.840 -4.770 ;
        RECT 92.300 -4.890 92.590 -4.770 ;
    END
  END WWLD[5]
  PIN WWLD[6]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 -7.630 4.730 -7.510 ;
        RECT 10.190 -7.630 10.480 -7.510 ;
        RECT 15.940 -7.630 16.230 -7.510 ;
        RECT 21.690 -7.630 21.980 -7.510 ;
        RECT 27.440 -7.630 27.730 -7.510 ;
        RECT 33.190 -7.630 33.480 -7.510 ;
        RECT 38.940 -7.630 39.230 -7.510 ;
        RECT 44.690 -7.630 44.980 -7.510 ;
        RECT 50.440 -7.630 50.730 -7.510 ;
        RECT 56.190 -7.630 56.480 -7.510 ;
        RECT 61.940 -7.630 62.230 -7.510 ;
        RECT 67.690 -7.630 67.980 -7.510 ;
        RECT 73.440 -7.630 73.730 -7.510 ;
        RECT 79.190 -7.630 79.480 -7.510 ;
        RECT 84.940 -7.630 85.230 -7.510 ;
        RECT 90.690 -7.630 90.980 -7.510 ;
        RECT -45.490 -7.770 94.660 -7.630 ;
        RECT 6.050 -7.890 6.340 -7.770 ;
        RECT 11.800 -7.890 12.090 -7.770 ;
        RECT 17.550 -7.890 17.840 -7.770 ;
        RECT 23.300 -7.890 23.590 -7.770 ;
        RECT 29.050 -7.890 29.340 -7.770 ;
        RECT 34.800 -7.890 35.090 -7.770 ;
        RECT 40.550 -7.890 40.840 -7.770 ;
        RECT 46.300 -7.890 46.590 -7.770 ;
        RECT 52.050 -7.890 52.340 -7.770 ;
        RECT 57.800 -7.890 58.090 -7.770 ;
        RECT 63.550 -7.890 63.840 -7.770 ;
        RECT 69.300 -7.890 69.590 -7.770 ;
        RECT 75.050 -7.890 75.340 -7.770 ;
        RECT 80.800 -7.890 81.090 -7.770 ;
        RECT 86.550 -7.890 86.840 -7.770 ;
        RECT 92.300 -7.890 92.590 -7.770 ;
    END
  END WWLD[6]
  PIN WWLD[7]
    ANTENNAGATEAREA 2.016000 ;
    PORT
      LAYER met1 ;
        RECT 4.440 -10.040 4.730 -9.920 ;
        RECT 10.190 -10.040 10.480 -9.920 ;
        RECT 15.940 -10.040 16.230 -9.920 ;
        RECT 21.690 -10.040 21.980 -9.920 ;
        RECT 27.440 -10.040 27.730 -9.920 ;
        RECT 33.190 -10.040 33.480 -9.920 ;
        RECT 38.940 -10.040 39.230 -9.920 ;
        RECT 44.690 -10.040 44.980 -9.920 ;
        RECT 50.440 -10.040 50.730 -9.920 ;
        RECT 56.190 -10.040 56.480 -9.920 ;
        RECT 61.940 -10.040 62.230 -9.920 ;
        RECT 67.690 -10.040 67.980 -9.920 ;
        RECT 73.440 -10.040 73.730 -9.920 ;
        RECT 79.190 -10.040 79.480 -9.920 ;
        RECT 84.940 -10.040 85.230 -9.920 ;
        RECT 90.690 -10.040 90.980 -9.920 ;
        RECT -45.490 -10.180 94.660 -10.040 ;
        RECT 6.050 -10.300 6.340 -10.180 ;
        RECT 11.800 -10.300 12.090 -10.180 ;
        RECT 17.550 -10.300 17.840 -10.180 ;
        RECT 23.300 -10.300 23.590 -10.180 ;
        RECT 29.050 -10.300 29.340 -10.180 ;
        RECT 34.800 -10.300 35.090 -10.180 ;
        RECT 40.550 -10.300 40.840 -10.180 ;
        RECT 46.300 -10.300 46.590 -10.180 ;
        RECT 52.050 -10.300 52.340 -10.180 ;
        RECT 57.800 -10.300 58.090 -10.180 ;
        RECT 63.550 -10.300 63.840 -10.180 ;
        RECT 69.300 -10.300 69.590 -10.180 ;
        RECT 75.050 -10.300 75.340 -10.180 ;
        RECT 80.800 -10.300 81.090 -10.180 ;
        RECT 86.550 -10.300 86.840 -10.180 ;
        RECT 92.300 -10.300 92.590 -10.180 ;
    END
  END WWLD[7]
  PIN SA_OUT[0]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 5.930 -6.070 6.290 -6.040 ;
        RECT 5.930 -6.370 100.480 -6.070 ;
        RECT 5.930 -6.400 6.290 -6.370 ;
    END
  END SA_OUT[0]
  PIN SA_OUT[1]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 11.680 -7.340 12.040 -7.310 ;
        RECT 11.680 -7.640 100.480 -7.340 ;
        RECT 11.680 -7.670 12.040 -7.640 ;
    END
  END SA_OUT[1]
  PIN SA_OUT[2]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 17.480 -8.710 17.840 -8.680 ;
        RECT 17.480 -9.010 100.480 -8.710 ;
        RECT 17.480 -9.040 17.840 -9.010 ;
    END
  END SA_OUT[2]
  PIN SA_OUT[3]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 23.180 -9.880 23.540 -9.850 ;
        RECT 23.180 -10.180 100.480 -9.880 ;
        RECT 23.180 -10.210 23.540 -10.180 ;
    END
  END SA_OUT[3]
  PIN SA_OUT[4]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 28.930 -11.130 29.290 -11.100 ;
        RECT 28.930 -11.430 100.480 -11.130 ;
        RECT 28.930 -11.460 29.290 -11.430 ;
    END
  END SA_OUT[4]
  PIN SA_OUT[5]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 34.680 -12.580 35.040 -12.550 ;
        RECT 34.680 -12.880 100.480 -12.580 ;
        RECT 34.680 -12.910 35.040 -12.880 ;
    END
  END SA_OUT[5]
  PIN SA_OUT[6]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 40.400 -13.800 40.800 -13.750 ;
        RECT 40.400 -14.100 100.480 -13.800 ;
        RECT 40.400 -14.150 40.800 -14.100 ;
    END
  END SA_OUT[6]
  PIN SA_OUT[7]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 46.180 -14.680 46.540 -14.650 ;
        RECT 46.180 -14.980 100.480 -14.680 ;
        RECT 46.180 -15.010 46.540 -14.980 ;
    END
  END SA_OUT[7]
  PIN SA_OUT[8]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 51.930 -15.510 52.290 -15.480 ;
        RECT 51.930 -15.810 100.480 -15.510 ;
        RECT 51.930 -15.840 52.290 -15.810 ;
    END
  END SA_OUT[8]
  PIN SA_OUT[9]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 57.680 -16.290 58.040 -16.260 ;
        RECT 57.680 -16.590 100.480 -16.290 ;
        RECT 57.680 -16.620 58.040 -16.590 ;
    END
  END SA_OUT[9]
  PIN SA_OUT[10]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 63.430 -17.150 63.790 -17.120 ;
        RECT 63.430 -17.450 100.480 -17.150 ;
        RECT 63.430 -17.480 63.790 -17.450 ;
    END
  END SA_OUT[10]
  PIN SA_OUT[11]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 69.180 -17.950 69.540 -17.920 ;
        RECT 69.180 -18.250 100.480 -17.950 ;
        RECT 69.180 -18.280 69.540 -18.250 ;
    END
  END SA_OUT[11]
  PIN SA_OUT[12]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 74.930 -18.750 75.290 -18.720 ;
        RECT 74.930 -19.050 100.480 -18.750 ;
        RECT 74.930 -19.080 75.290 -19.050 ;
    END
  END SA_OUT[12]
  PIN SA_OUT[13]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 80.680 -19.400 81.040 -19.370 ;
        RECT 80.680 -19.700 100.480 -19.400 ;
        RECT 80.680 -19.730 81.040 -19.700 ;
    END
  END SA_OUT[13]
  PIN SA_OUT[14]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 86.430 -20.540 86.790 -20.510 ;
        RECT 86.430 -20.840 100.480 -20.540 ;
        RECT 86.430 -20.870 86.790 -20.840 ;
    END
  END SA_OUT[14]
  PIN SA_OUT[15]
    ANTENNAGATEAREA 0.750000 ;
    ANTENNADIFFAREA 1.890000 ;
    PORT
      LAYER met3 ;
        RECT 92.180 -21.430 92.540 -21.400 ;
        RECT 92.180 -21.730 100.480 -21.430 ;
        RECT 92.180 -21.760 92.540 -21.730 ;
    END
  END SA_OUT[15]
  PIN EN
    ANTENNAGATEAREA 1.536000 ;
    PORT
      LAYER met3 ;
        RECT 7.300 -24.190 7.700 -24.140 ;
        RECT 8.850 -24.190 9.250 -24.140 ;
        RECT 18.800 -24.190 19.200 -24.140 ;
        RECT 20.350 -24.190 20.750 -24.140 ;
        RECT 30.300 -24.190 30.700 -24.140 ;
        RECT 31.840 -24.190 32.240 -24.140 ;
        RECT 41.770 -24.190 42.170 -24.140 ;
        RECT 43.360 -24.190 43.760 -24.150 ;
        RECT 53.290 -24.190 53.690 -24.140 ;
        RECT 54.840 -24.190 55.240 -24.140 ;
        RECT 64.800 -24.190 65.200 -24.150 ;
        RECT 66.330 -24.190 66.730 -24.150 ;
        RECT 76.310 -24.190 76.710 -24.140 ;
        RECT 77.840 -24.190 78.240 -24.140 ;
        RECT 87.800 -24.190 88.200 -24.140 ;
        RECT 89.320 -24.190 89.720 -24.130 ;
        RECT -45.420 -24.490 89.720 -24.190 ;
        RECT 7.300 -24.540 7.700 -24.490 ;
        RECT 8.850 -24.540 9.250 -24.490 ;
        RECT 18.800 -24.540 19.200 -24.490 ;
        RECT 20.350 -24.540 20.750 -24.490 ;
        RECT 30.300 -24.540 30.700 -24.490 ;
        RECT 31.840 -24.540 32.240 -24.490 ;
        RECT 41.770 -24.540 42.170 -24.490 ;
        RECT 43.360 -24.550 43.760 -24.490 ;
        RECT 53.290 -24.540 53.690 -24.490 ;
        RECT 54.840 -24.540 55.240 -24.490 ;
        RECT 64.800 -24.550 65.200 -24.490 ;
        RECT 66.330 -24.550 66.730 -24.490 ;
        RECT 76.310 -24.540 76.710 -24.490 ;
        RECT 77.840 -24.540 78.240 -24.490 ;
        RECT 87.800 -24.540 88.200 -24.490 ;
        RECT 89.320 -24.540 89.720 -24.490 ;
    END
  END EN
  PIN PRE_A
    ANTENNAGATEAREA 1.008000 ;
    PORT
      LAYER met3 ;
        RECT 4.610 -24.950 5.010 -24.910 ;
        RECT 11.540 -24.950 11.940 -24.840 ;
        RECT 16.100 -24.950 16.500 -24.830 ;
        RECT 23.030 -24.950 23.430 -24.880 ;
        RECT 27.620 -24.950 28.020 -24.890 ;
        RECT 34.540 -24.950 34.940 -24.870 ;
        RECT 39.120 -24.950 39.520 -24.890 ;
        RECT 46.030 -24.950 46.430 -24.910 ;
        RECT 50.610 -24.950 51.010 -24.850 ;
        RECT 57.540 -24.950 57.940 -24.870 ;
        RECT 62.110 -24.950 62.510 -24.830 ;
        RECT 69.030 -24.950 69.430 -24.870 ;
        RECT 73.610 -24.950 74.010 -24.870 ;
        RECT 80.530 -24.950 80.930 -24.900 ;
        RECT 85.110 -24.950 85.510 -24.890 ;
        RECT 92.030 -24.950 92.390 -24.870 ;
        RECT -45.420 -25.250 92.390 -24.950 ;
        RECT 4.610 -25.310 5.010 -25.250 ;
        RECT 23.030 -25.280 23.430 -25.250 ;
        RECT 27.620 -25.290 28.020 -25.250 ;
        RECT 34.540 -25.270 34.940 -25.250 ;
        RECT 39.120 -25.290 39.520 -25.250 ;
        RECT 46.030 -25.310 46.430 -25.250 ;
        RECT 57.540 -25.270 57.940 -25.250 ;
        RECT 69.030 -25.270 69.430 -25.250 ;
        RECT 73.610 -25.270 74.010 -25.250 ;
        RECT 80.530 -25.300 80.930 -25.250 ;
        RECT 85.110 -25.290 85.510 -25.250 ;
    END
  END PRE_A
  PIN VDD
    ANTENNADIFFAREA 415.516785 ;
    PORT
      LAYER nwell ;
        RECT 2.250 48.670 94.660 50.590 ;
        RECT 4.700 -11.420 6.080 48.670 ;
        RECT 10.450 -11.420 11.830 48.670 ;
        RECT 16.200 -11.420 17.580 48.670 ;
        RECT 21.950 -11.420 23.330 48.670 ;
        RECT 27.700 -11.420 29.080 48.670 ;
        RECT 33.450 -11.420 34.830 48.670 ;
        RECT 39.200 -11.420 40.580 48.670 ;
        RECT 44.950 -11.420 46.330 48.670 ;
        RECT 50.700 -11.420 52.080 48.670 ;
        RECT 56.450 -11.420 57.830 48.670 ;
        RECT 62.200 -11.420 63.580 48.670 ;
        RECT 67.950 -11.420 69.330 48.670 ;
        RECT 73.700 -11.420 75.080 48.670 ;
        RECT 79.450 -11.420 80.830 48.670 ;
        RECT 85.200 -11.420 86.580 48.670 ;
        RECT 90.950 -11.420 92.330 48.670 ;
        RECT 2.250 -14.140 94.660 -11.420 ;
        RECT 2.250 -22.560 94.660 -21.210 ;
        RECT 2.250 -24.540 5.890 -22.560 ;
        RECT 10.640 -24.540 17.390 -22.560 ;
        RECT 22.140 -24.540 28.890 -22.560 ;
        RECT 33.640 -24.540 40.390 -22.560 ;
        RECT 45.140 -24.540 51.890 -22.560 ;
        RECT 56.640 -24.540 63.390 -22.560 ;
        RECT 68.140 -24.540 74.890 -22.560 ;
        RECT 79.640 -24.540 86.390 -22.560 ;
        RECT 91.140 -24.540 94.660 -22.560 ;
        RECT -38.440 -36.140 -31.820 -31.170 ;
        RECT -26.940 -36.140 -20.320 -31.170 ;
        RECT -3.310 -36.140 3.310 -31.170 ;
        RECT 8.500 -36.140 15.120 -31.170 ;
        RECT 20.320 -36.140 26.940 -31.170 ;
        RECT 32.140 -36.140 38.760 -31.170 ;
        RECT 43.960 -36.140 50.580 -31.170 ;
        RECT 55.780 -36.140 62.400 -31.170 ;
        RECT 67.600 -36.140 74.220 -31.170 ;
        RECT 79.420 -36.140 86.040 -31.170 ;
        RECT 91.260 -36.140 97.880 -31.170 ;
        RECT 103.100 -36.140 109.720 -31.170 ;
        RECT 114.970 -36.140 121.590 -31.170 ;
        RECT 126.840 -36.140 133.460 -31.170 ;
        RECT 135.850 -36.140 142.470 -31.170 ;
        RECT -38.440 -63.470 -31.820 -53.940 ;
        RECT -26.940 -63.470 -20.320 -53.940 ;
        RECT -3.310 -63.470 3.310 -53.940 ;
        RECT 8.500 -63.470 15.120 -53.940 ;
        RECT 20.320 -63.470 26.940 -53.940 ;
        RECT 32.140 -63.470 38.760 -53.940 ;
        RECT 43.960 -63.470 50.580 -53.940 ;
        RECT 55.780 -63.470 62.400 -53.940 ;
        RECT 67.600 -63.470 74.220 -53.940 ;
        RECT 79.420 -63.470 86.040 -53.940 ;
        RECT 91.260 -63.470 97.880 -53.940 ;
        RECT 103.100 -63.470 109.720 -53.940 ;
        RECT 114.970 -63.470 121.590 -53.940 ;
        RECT 126.840 -63.470 133.460 -53.940 ;
        RECT 135.850 -63.470 142.470 -53.940 ;
        RECT -38.440 -86.240 -31.820 -81.270 ;
        RECT -26.940 -86.240 -20.320 -81.270 ;
        RECT -3.310 -86.240 3.310 -81.270 ;
        RECT 8.500 -86.240 15.120 -81.270 ;
        RECT 20.320 -86.240 26.940 -81.270 ;
        RECT 32.140 -86.240 38.760 -81.270 ;
        RECT 43.960 -86.240 50.580 -81.270 ;
        RECT 55.780 -86.240 62.400 -81.270 ;
        RECT 67.600 -86.240 74.220 -81.270 ;
        RECT 79.420 -86.240 86.040 -81.270 ;
        RECT 91.260 -86.240 97.880 -81.270 ;
        RECT 103.100 -86.240 109.720 -81.270 ;
        RECT 114.970 -86.240 121.590 -81.270 ;
        RECT 126.840 -86.240 133.460 -81.270 ;
        RECT 135.850 -86.240 142.470 -81.270 ;
      LAYER met3 ;
        RECT 5.190 50.640 5.590 50.740 ;
        RECT 10.950 50.640 11.350 50.740 ;
        RECT 16.700 50.640 17.100 50.740 ;
        RECT 22.430 50.640 22.830 50.740 ;
        RECT 28.190 50.640 28.590 50.740 ;
        RECT 33.930 50.640 34.330 50.740 ;
        RECT 39.680 50.640 40.080 50.740 ;
        RECT 45.430 50.640 45.830 50.740 ;
        RECT 51.180 50.640 51.580 50.740 ;
        RECT 56.940 50.640 57.340 50.740 ;
        RECT 62.690 50.640 63.090 50.730 ;
        RECT 68.430 50.640 68.830 50.740 ;
        RECT 74.180 50.640 74.580 50.740 ;
        RECT 79.930 50.640 80.330 50.740 ;
        RECT 85.670 50.640 86.070 50.740 ;
        RECT 91.420 50.640 91.820 50.740 ;
        RECT -45.490 50.340 100.380 50.640 ;
        RECT -43.170 50.280 -42.810 50.340 ;
        RECT 62.690 50.330 63.090 50.340 ;
        RECT -43.170 -30.670 -42.810 -30.600 ;
        RECT -35.270 -30.670 -34.910 -30.640 ;
        RECT -23.770 -30.670 -23.410 -30.640 ;
        RECT 11.670 -30.670 12.030 -30.660 ;
        RECT 47.130 -30.670 47.490 -30.640 ;
        RECT 82.590 -30.670 82.950 -30.650 ;
        RECT 94.430 -30.670 94.790 -30.660 ;
        RECT 118.140 -30.670 118.500 -30.630 ;
        RECT 130.010 -30.670 130.370 -30.650 ;
        RECT -45.150 -30.970 144.360 -30.670 ;
        RECT -35.270 -31.000 -34.910 -30.970 ;
        RECT -23.770 -31.000 -23.410 -30.970 ;
        RECT -0.140 -31.040 0.220 -30.970 ;
        RECT 11.670 -31.020 12.030 -30.970 ;
        RECT 23.490 -31.030 23.850 -30.970 ;
        RECT 35.310 -31.030 35.670 -30.970 ;
        RECT 47.130 -31.000 47.490 -30.970 ;
        RECT 58.950 -31.030 59.310 -30.970 ;
        RECT 70.770 -31.030 71.130 -30.970 ;
        RECT 82.590 -31.010 82.950 -30.970 ;
        RECT 94.430 -31.020 94.790 -30.970 ;
        RECT 106.270 -31.030 106.630 -30.970 ;
        RECT 118.140 -30.990 118.500 -30.970 ;
        RECT 130.010 -31.010 130.370 -30.970 ;
        RECT 139.020 -31.030 139.380 -30.970 ;
    END
  END VDD
  PIN VSS
    ANTENNAGATEAREA 16.128000 ;
    ANTENNADIFFAREA 316.692780 ;
    PORT
      LAYER pwell ;
        RECT 2.250 33.560 4.700 48.670 ;
        RECT 2.240 33.420 4.700 33.560 ;
        RECT 2.250 28.740 4.700 33.420 ;
        RECT 2.240 28.600 4.700 28.740 ;
        RECT 2.250 -11.420 4.700 28.600 ;
        RECT 6.080 -11.420 10.450 48.670 ;
        RECT 11.830 -11.420 16.200 48.670 ;
        RECT 17.580 -11.420 21.950 48.670 ;
        RECT 23.330 -11.420 27.700 48.670 ;
        RECT 29.080 -11.420 33.450 48.670 ;
        RECT 34.830 -11.420 39.200 48.670 ;
        RECT 40.580 -11.420 44.950 48.670 ;
        RECT 46.330 -11.420 50.700 48.670 ;
        RECT 52.080 -11.420 56.450 48.670 ;
        RECT 57.830 -11.420 62.200 48.670 ;
        RECT 63.580 -11.420 67.950 48.670 ;
        RECT 69.330 -11.420 73.700 48.670 ;
        RECT 75.080 -11.420 79.450 48.670 ;
        RECT 80.830 -11.420 85.200 48.670 ;
        RECT 86.580 -11.420 90.950 48.670 ;
        RECT 92.330 -11.420 94.660 48.670 ;
        RECT 2.250 -21.210 94.660 -14.140 ;
        RECT 5.890 -24.540 10.640 -22.560 ;
        RECT 17.390 -24.540 22.140 -22.560 ;
        RECT 28.890 -24.540 33.640 -22.560 ;
        RECT 40.390 -24.540 45.140 -22.560 ;
        RECT 51.890 -24.540 56.640 -22.560 ;
        RECT 63.390 -24.540 68.140 -22.560 ;
        RECT 74.890 -24.540 79.640 -22.560 ;
        RECT 86.390 -24.540 91.140 -22.560 ;
        RECT -38.440 -53.940 -31.820 -36.140 ;
        RECT -26.940 -53.940 -20.320 -36.140 ;
        RECT -15.120 -53.940 -8.500 -36.140 ;
        RECT -3.310 -53.940 3.310 -36.140 ;
        RECT 8.500 -53.940 15.120 -36.140 ;
        RECT 20.320 -53.940 26.940 -36.140 ;
        RECT 32.140 -53.940 38.760 -36.140 ;
        RECT 43.960 -53.940 50.580 -36.140 ;
        RECT 55.780 -53.940 62.400 -36.140 ;
        RECT 67.600 -53.940 74.220 -36.140 ;
        RECT 79.420 -53.940 86.040 -36.140 ;
        RECT 91.260 -53.940 97.880 -36.140 ;
        RECT 103.100 -53.940 109.720 -36.140 ;
        RECT 114.970 -53.940 121.590 -36.140 ;
        RECT 126.840 -53.940 133.460 -36.140 ;
        RECT 135.850 -53.940 142.470 -36.140 ;
        RECT -38.440 -81.270 -31.820 -63.470 ;
        RECT -26.940 -81.270 -20.320 -63.470 ;
        RECT -15.120 -81.270 -8.500 -63.470 ;
        RECT -3.310 -81.270 3.310 -63.470 ;
        RECT 8.500 -81.270 15.120 -63.470 ;
        RECT 20.320 -81.270 26.940 -63.470 ;
        RECT 32.140 -81.270 38.760 -63.470 ;
        RECT 43.960 -81.270 50.580 -63.470 ;
        RECT 55.780 -81.270 62.400 -63.470 ;
        RECT 67.600 -81.270 74.220 -63.470 ;
        RECT 79.420 -81.270 86.040 -63.470 ;
        RECT 91.260 -81.270 97.880 -63.470 ;
        RECT 103.100 -81.270 109.720 -63.470 ;
        RECT 114.970 -81.270 121.590 -63.470 ;
        RECT 126.840 -81.270 133.460 -63.470 ;
        RECT 135.850 -81.270 142.470 -63.470 ;
      LAYER met3 ;
        RECT -0.400 -20.300 0.000 -20.250 ;
        RECT -45.520 -20.600 0.000 -20.300 ;
        RECT -41.830 -20.670 -41.470 -20.600 ;
        RECT -0.400 -20.650 0.000 -20.600 ;
        RECT -0.350 -23.210 -0.050 -20.650 ;
        RECT 8.060 -23.200 8.460 -23.150 ;
        RECT 8.050 -23.210 8.460 -23.200 ;
        RECT 19.550 -23.210 19.950 -23.160 ;
        RECT 30.980 -23.210 31.380 -23.170 ;
        RECT 42.550 -23.210 42.950 -23.180 ;
        RECT 53.950 -23.210 54.350 -23.160 ;
        RECT 65.630 -23.210 66.030 -23.160 ;
        RECT 77.080 -23.210 77.480 -23.160 ;
        RECT 88.650 -23.190 89.050 -23.140 ;
        RECT 88.640 -23.210 89.050 -23.190 ;
        RECT -0.350 -23.510 89.050 -23.210 ;
        RECT 8.060 -23.550 8.460 -23.510 ;
        RECT 19.550 -23.560 19.950 -23.510 ;
        RECT 30.970 -23.520 31.380 -23.510 ;
        RECT 30.980 -23.570 31.380 -23.520 ;
        RECT 42.540 -23.530 42.950 -23.510 ;
        RECT 42.550 -23.580 42.950 -23.530 ;
        RECT 53.950 -23.560 54.350 -23.510 ;
        RECT 65.630 -23.560 66.030 -23.510 ;
        RECT 77.080 -23.560 77.480 -23.510 ;
        RECT 88.650 -23.540 89.050 -23.510 ;
    END
  END VSS
  PIN Iref0
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER met2 ;
        RECT 144.460 -44.740 144.720 -44.420 ;
        RECT 144.510 -90.100 144.680 -44.740 ;
    END
  END Iref0
  PIN Iref1
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER met2 ;
        RECT 145.020 -45.630 145.280 -45.310 ;
        RECT 145.070 -90.100 145.240 -45.630 ;
    END
  END Iref1
  PIN Iref2
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER met2 ;
        RECT 145.560 -72.000 145.820 -71.680 ;
        RECT 145.610 -90.100 145.780 -72.000 ;
    END
  END Iref2
  PIN Iref3
    ANTENNAGATEAREA 16.000000 ;
    PORT
      LAYER met2 ;
        RECT 146.110 -72.970 146.370 -72.650 ;
        RECT 146.160 -90.100 146.330 -72.970 ;
    END
  END Iref3
  OBS
      LAYER nwell ;
        RECT -15.120 -36.140 -8.500 -31.170 ;
        RECT -15.120 -63.470 -8.500 -53.940 ;
        RECT -15.120 -86.240 -8.500 -81.270 ;
      LAYER li1 ;
        RECT 4.340 49.990 4.670 50.160 ;
        RECT 5.210 49.990 5.540 50.160 ;
        RECT 6.080 49.990 6.410 50.160 ;
        RECT 10.090 49.990 10.420 50.160 ;
        RECT 10.960 49.990 11.290 50.160 ;
        RECT 11.830 49.990 12.160 50.160 ;
        RECT 15.840 49.990 16.170 50.160 ;
        RECT 16.710 49.990 17.040 50.160 ;
        RECT 17.580 49.990 17.910 50.160 ;
        RECT 21.590 49.990 21.920 50.160 ;
        RECT 22.460 49.990 22.790 50.160 ;
        RECT 23.330 49.990 23.660 50.160 ;
        RECT 27.340 49.990 27.670 50.160 ;
        RECT 28.210 49.990 28.540 50.160 ;
        RECT 29.080 49.990 29.410 50.160 ;
        RECT 33.090 49.990 33.420 50.160 ;
        RECT 33.960 49.990 34.290 50.160 ;
        RECT 34.830 49.990 35.160 50.160 ;
        RECT 38.840 49.990 39.170 50.160 ;
        RECT 39.710 49.990 40.040 50.160 ;
        RECT 40.580 49.990 40.910 50.160 ;
        RECT 44.590 49.990 44.920 50.160 ;
        RECT 45.460 49.990 45.790 50.160 ;
        RECT 46.330 49.990 46.660 50.160 ;
        RECT 50.340 49.990 50.670 50.160 ;
        RECT 51.210 49.990 51.540 50.160 ;
        RECT 52.080 49.990 52.410 50.160 ;
        RECT 56.090 49.990 56.420 50.160 ;
        RECT 56.960 49.990 57.290 50.160 ;
        RECT 57.830 49.990 58.160 50.160 ;
        RECT 61.840 49.990 62.170 50.160 ;
        RECT 62.710 49.990 63.040 50.160 ;
        RECT 63.580 49.990 63.910 50.160 ;
        RECT 67.590 49.990 67.920 50.160 ;
        RECT 68.460 49.990 68.790 50.160 ;
        RECT 69.330 49.990 69.660 50.160 ;
        RECT 73.340 49.990 73.670 50.160 ;
        RECT 74.210 49.990 74.540 50.160 ;
        RECT 75.080 49.990 75.410 50.160 ;
        RECT 79.090 49.990 79.420 50.160 ;
        RECT 79.960 49.990 80.290 50.160 ;
        RECT 80.830 49.990 81.160 50.160 ;
        RECT 84.840 49.990 85.170 50.160 ;
        RECT 85.710 49.990 86.040 50.160 ;
        RECT 86.580 49.990 86.910 50.160 ;
        RECT 90.590 49.990 90.920 50.160 ;
        RECT 91.460 49.990 91.790 50.160 ;
        RECT 92.330 49.990 92.660 50.160 ;
        RECT 4.110 49.340 4.280 49.750 ;
        RECT 4.550 49.650 4.720 49.750 ;
        RECT 6.030 49.650 6.200 49.750 ;
        RECT 4.550 49.480 6.200 49.650 ;
        RECT 4.550 49.350 4.720 49.480 ;
        RECT 6.030 49.350 6.200 49.480 ;
        RECT 4.100 49.170 4.280 49.340 ;
        RECT 5.070 49.170 5.240 49.290 ;
        RECT 4.100 49.000 5.240 49.170 ;
        RECT 5.070 48.870 5.240 49.000 ;
        RECT 5.510 49.180 5.680 49.290 ;
        RECT 6.470 49.180 6.640 49.750 ;
        RECT 9.860 49.340 10.030 49.750 ;
        RECT 10.300 49.650 10.470 49.750 ;
        RECT 11.780 49.650 11.950 49.750 ;
        RECT 10.300 49.480 11.950 49.650 ;
        RECT 10.300 49.350 10.470 49.480 ;
        RECT 11.780 49.350 11.950 49.480 ;
        RECT 5.510 48.990 6.640 49.180 ;
        RECT 9.850 49.170 10.030 49.340 ;
        RECT 10.820 49.170 10.990 49.290 ;
        RECT 9.850 49.000 10.990 49.170 ;
        RECT 5.510 48.870 5.680 48.990 ;
        RECT 10.820 48.870 10.990 49.000 ;
        RECT 11.260 49.180 11.430 49.290 ;
        RECT 12.220 49.180 12.390 49.750 ;
        RECT 15.610 49.340 15.780 49.750 ;
        RECT 16.050 49.650 16.220 49.750 ;
        RECT 17.530 49.650 17.700 49.750 ;
        RECT 16.050 49.480 17.700 49.650 ;
        RECT 16.050 49.350 16.220 49.480 ;
        RECT 17.530 49.350 17.700 49.480 ;
        RECT 11.260 48.990 12.390 49.180 ;
        RECT 15.600 49.170 15.780 49.340 ;
        RECT 16.570 49.170 16.740 49.290 ;
        RECT 15.600 49.000 16.740 49.170 ;
        RECT 11.260 48.870 11.430 48.990 ;
        RECT 16.570 48.870 16.740 49.000 ;
        RECT 17.010 49.180 17.180 49.290 ;
        RECT 17.970 49.180 18.140 49.750 ;
        RECT 21.360 49.340 21.530 49.750 ;
        RECT 21.800 49.650 21.970 49.750 ;
        RECT 23.280 49.650 23.450 49.750 ;
        RECT 21.800 49.480 23.450 49.650 ;
        RECT 21.800 49.350 21.970 49.480 ;
        RECT 23.280 49.350 23.450 49.480 ;
        RECT 17.010 48.990 18.140 49.180 ;
        RECT 21.350 49.170 21.530 49.340 ;
        RECT 22.320 49.170 22.490 49.290 ;
        RECT 21.350 49.000 22.490 49.170 ;
        RECT 17.010 48.870 17.180 48.990 ;
        RECT 22.320 48.870 22.490 49.000 ;
        RECT 22.760 49.180 22.930 49.290 ;
        RECT 23.720 49.180 23.890 49.750 ;
        RECT 27.110 49.340 27.280 49.750 ;
        RECT 27.550 49.650 27.720 49.750 ;
        RECT 29.030 49.650 29.200 49.750 ;
        RECT 27.550 49.480 29.200 49.650 ;
        RECT 27.550 49.350 27.720 49.480 ;
        RECT 29.030 49.350 29.200 49.480 ;
        RECT 22.760 48.990 23.890 49.180 ;
        RECT 27.100 49.170 27.280 49.340 ;
        RECT 28.070 49.170 28.240 49.290 ;
        RECT 27.100 49.000 28.240 49.170 ;
        RECT 22.760 48.870 22.930 48.990 ;
        RECT 28.070 48.870 28.240 49.000 ;
        RECT 28.510 49.180 28.680 49.290 ;
        RECT 29.470 49.180 29.640 49.750 ;
        RECT 32.860 49.340 33.030 49.750 ;
        RECT 33.300 49.650 33.470 49.750 ;
        RECT 34.780 49.650 34.950 49.750 ;
        RECT 33.300 49.480 34.950 49.650 ;
        RECT 33.300 49.350 33.470 49.480 ;
        RECT 34.780 49.350 34.950 49.480 ;
        RECT 28.510 48.990 29.640 49.180 ;
        RECT 32.850 49.170 33.030 49.340 ;
        RECT 33.820 49.170 33.990 49.290 ;
        RECT 32.850 49.000 33.990 49.170 ;
        RECT 28.510 48.870 28.680 48.990 ;
        RECT 33.820 48.870 33.990 49.000 ;
        RECT 34.260 49.180 34.430 49.290 ;
        RECT 35.220 49.180 35.390 49.750 ;
        RECT 38.610 49.340 38.780 49.750 ;
        RECT 39.050 49.650 39.220 49.750 ;
        RECT 40.530 49.650 40.700 49.750 ;
        RECT 39.050 49.480 40.700 49.650 ;
        RECT 39.050 49.350 39.220 49.480 ;
        RECT 40.530 49.350 40.700 49.480 ;
        RECT 34.260 48.990 35.390 49.180 ;
        RECT 38.600 49.170 38.780 49.340 ;
        RECT 39.570 49.170 39.740 49.290 ;
        RECT 38.600 49.000 39.740 49.170 ;
        RECT 34.260 48.870 34.430 48.990 ;
        RECT 39.570 48.870 39.740 49.000 ;
        RECT 40.010 49.180 40.180 49.290 ;
        RECT 40.970 49.180 41.140 49.750 ;
        RECT 44.360 49.340 44.530 49.750 ;
        RECT 44.800 49.650 44.970 49.750 ;
        RECT 46.280 49.650 46.450 49.750 ;
        RECT 44.800 49.480 46.450 49.650 ;
        RECT 44.800 49.350 44.970 49.480 ;
        RECT 46.280 49.350 46.450 49.480 ;
        RECT 40.010 48.990 41.140 49.180 ;
        RECT 44.350 49.170 44.530 49.340 ;
        RECT 45.320 49.170 45.490 49.290 ;
        RECT 44.350 49.000 45.490 49.170 ;
        RECT 40.010 48.870 40.180 48.990 ;
        RECT 45.320 48.870 45.490 49.000 ;
        RECT 45.760 49.180 45.930 49.290 ;
        RECT 46.720 49.180 46.890 49.750 ;
        RECT 50.110 49.340 50.280 49.750 ;
        RECT 50.550 49.650 50.720 49.750 ;
        RECT 52.030 49.650 52.200 49.750 ;
        RECT 50.550 49.480 52.200 49.650 ;
        RECT 50.550 49.350 50.720 49.480 ;
        RECT 52.030 49.350 52.200 49.480 ;
        RECT 45.760 48.990 46.890 49.180 ;
        RECT 50.100 49.170 50.280 49.340 ;
        RECT 51.070 49.170 51.240 49.290 ;
        RECT 50.100 49.000 51.240 49.170 ;
        RECT 45.760 48.870 45.930 48.990 ;
        RECT 51.070 48.870 51.240 49.000 ;
        RECT 51.510 49.180 51.680 49.290 ;
        RECT 52.470 49.180 52.640 49.750 ;
        RECT 55.860 49.340 56.030 49.750 ;
        RECT 56.300 49.650 56.470 49.750 ;
        RECT 57.780 49.650 57.950 49.750 ;
        RECT 56.300 49.480 57.950 49.650 ;
        RECT 56.300 49.350 56.470 49.480 ;
        RECT 57.780 49.350 57.950 49.480 ;
        RECT 51.510 48.990 52.640 49.180 ;
        RECT 55.850 49.170 56.030 49.340 ;
        RECT 56.820 49.170 56.990 49.290 ;
        RECT 55.850 49.000 56.990 49.170 ;
        RECT 51.510 48.870 51.680 48.990 ;
        RECT 56.820 48.870 56.990 49.000 ;
        RECT 57.260 49.180 57.430 49.290 ;
        RECT 58.220 49.180 58.390 49.750 ;
        RECT 61.610 49.340 61.780 49.750 ;
        RECT 62.050 49.650 62.220 49.750 ;
        RECT 63.530 49.650 63.700 49.750 ;
        RECT 62.050 49.480 63.700 49.650 ;
        RECT 62.050 49.350 62.220 49.480 ;
        RECT 63.530 49.350 63.700 49.480 ;
        RECT 57.260 48.990 58.390 49.180 ;
        RECT 61.600 49.170 61.780 49.340 ;
        RECT 62.570 49.170 62.740 49.290 ;
        RECT 61.600 49.000 62.740 49.170 ;
        RECT 57.260 48.870 57.430 48.990 ;
        RECT 62.570 48.870 62.740 49.000 ;
        RECT 63.010 49.180 63.180 49.290 ;
        RECT 63.970 49.180 64.140 49.750 ;
        RECT 67.360 49.340 67.530 49.750 ;
        RECT 67.800 49.650 67.970 49.750 ;
        RECT 69.280 49.650 69.450 49.750 ;
        RECT 67.800 49.480 69.450 49.650 ;
        RECT 67.800 49.350 67.970 49.480 ;
        RECT 69.280 49.350 69.450 49.480 ;
        RECT 63.010 48.990 64.140 49.180 ;
        RECT 67.350 49.170 67.530 49.340 ;
        RECT 68.320 49.170 68.490 49.290 ;
        RECT 67.350 49.000 68.490 49.170 ;
        RECT 63.010 48.870 63.180 48.990 ;
        RECT 68.320 48.870 68.490 49.000 ;
        RECT 68.760 49.180 68.930 49.290 ;
        RECT 69.720 49.180 69.890 49.750 ;
        RECT 73.110 49.340 73.280 49.750 ;
        RECT 73.550 49.650 73.720 49.750 ;
        RECT 75.030 49.650 75.200 49.750 ;
        RECT 73.550 49.480 75.200 49.650 ;
        RECT 73.550 49.350 73.720 49.480 ;
        RECT 75.030 49.350 75.200 49.480 ;
        RECT 68.760 48.990 69.890 49.180 ;
        RECT 73.100 49.170 73.280 49.340 ;
        RECT 74.070 49.170 74.240 49.290 ;
        RECT 73.100 49.000 74.240 49.170 ;
        RECT 68.760 48.870 68.930 48.990 ;
        RECT 74.070 48.870 74.240 49.000 ;
        RECT 74.510 49.180 74.680 49.290 ;
        RECT 75.470 49.180 75.640 49.750 ;
        RECT 78.860 49.340 79.030 49.750 ;
        RECT 79.300 49.650 79.470 49.750 ;
        RECT 80.780 49.650 80.950 49.750 ;
        RECT 79.300 49.480 80.950 49.650 ;
        RECT 79.300 49.350 79.470 49.480 ;
        RECT 80.780 49.350 80.950 49.480 ;
        RECT 74.510 48.990 75.640 49.180 ;
        RECT 78.850 49.170 79.030 49.340 ;
        RECT 79.820 49.170 79.990 49.290 ;
        RECT 78.850 49.000 79.990 49.170 ;
        RECT 74.510 48.870 74.680 48.990 ;
        RECT 79.820 48.870 79.990 49.000 ;
        RECT 80.260 49.180 80.430 49.290 ;
        RECT 81.220 49.180 81.390 49.750 ;
        RECT 84.610 49.340 84.780 49.750 ;
        RECT 85.050 49.650 85.220 49.750 ;
        RECT 86.530 49.650 86.700 49.750 ;
        RECT 85.050 49.480 86.700 49.650 ;
        RECT 85.050 49.350 85.220 49.480 ;
        RECT 86.530 49.350 86.700 49.480 ;
        RECT 80.260 48.990 81.390 49.180 ;
        RECT 84.600 49.170 84.780 49.340 ;
        RECT 85.570 49.170 85.740 49.290 ;
        RECT 84.600 49.000 85.740 49.170 ;
        RECT 80.260 48.870 80.430 48.990 ;
        RECT 85.570 48.870 85.740 49.000 ;
        RECT 86.010 49.180 86.180 49.290 ;
        RECT 86.970 49.180 87.140 49.750 ;
        RECT 90.360 49.340 90.530 49.750 ;
        RECT 90.800 49.650 90.970 49.750 ;
        RECT 92.280 49.650 92.450 49.750 ;
        RECT 90.800 49.480 92.450 49.650 ;
        RECT 90.800 49.350 90.970 49.480 ;
        RECT 92.280 49.350 92.450 49.480 ;
        RECT 86.010 48.990 87.140 49.180 ;
        RECT 90.350 49.170 90.530 49.340 ;
        RECT 91.320 49.170 91.490 49.290 ;
        RECT 90.350 49.000 91.490 49.170 ;
        RECT 86.010 48.870 86.180 48.990 ;
        RECT 91.320 48.870 91.490 49.000 ;
        RECT 91.760 49.180 91.930 49.290 ;
        RECT 92.720 49.180 92.890 49.750 ;
        RECT 91.760 48.990 92.890 49.180 ;
        RECT 91.760 48.870 91.930 48.990 ;
        RECT 2.990 48.130 3.250 48.220 ;
        RECT 3.900 48.130 4.160 48.220 ;
        RECT 2.900 47.920 3.320 48.130 ;
        RECT 3.830 47.920 4.250 48.130 ;
        RECT 2.520 47.530 2.690 47.860 ;
        RECT 4.500 47.260 4.670 47.950 ;
        RECT 5.040 47.090 5.210 47.960 ;
        RECT 5.480 47.920 5.900 48.200 ;
        RECT 7.120 48.090 7.290 48.420 ;
        RECT 8.740 48.130 9.000 48.220 ;
        RECT 9.650 48.130 9.910 48.220 ;
        RECT 6.420 47.920 7.840 48.090 ;
        RECT 8.650 47.920 9.070 48.130 ;
        RECT 9.580 47.920 10.000 48.130 ;
        RECT 5.480 47.480 7.060 47.650 ;
        RECT 8.270 47.530 8.440 47.860 ;
        RECT 3.720 46.920 5.300 47.090 ;
        RECT 2.900 46.480 4.360 46.650 ;
        RECT 3.360 46.420 3.650 46.480 ;
        RECT 4.880 46.310 5.300 46.650 ;
        RECT 5.560 46.610 5.730 47.480 ;
        RECT 6.110 46.610 6.280 47.300 ;
        RECT 10.250 47.260 10.420 47.950 ;
        RECT 10.790 47.090 10.960 47.960 ;
        RECT 11.230 47.920 11.650 48.200 ;
        RECT 12.870 48.090 13.040 48.420 ;
        RECT 14.490 48.130 14.750 48.220 ;
        RECT 15.400 48.130 15.660 48.220 ;
        RECT 12.170 47.920 13.590 48.090 ;
        RECT 14.400 47.920 14.820 48.130 ;
        RECT 15.330 47.920 15.750 48.130 ;
        RECT 11.230 47.480 12.810 47.650 ;
        RECT 14.020 47.530 14.190 47.860 ;
        RECT 8.060 46.710 8.230 47.040 ;
        RECT 9.470 46.920 11.050 47.090 ;
        RECT 6.530 46.440 6.950 46.650 ;
        RECT 7.420 46.440 7.840 46.650 ;
        RECT 8.650 46.480 10.110 46.650 ;
        RECT 6.600 46.380 6.860 46.440 ;
        RECT 7.510 46.380 7.770 46.440 ;
        RECT 9.110 46.420 9.400 46.480 ;
        RECT 10.630 46.310 11.050 46.650 ;
        RECT 11.310 46.610 11.480 47.480 ;
        RECT 11.860 46.610 12.030 47.300 ;
        RECT 16.000 47.260 16.170 47.950 ;
        RECT 16.540 47.090 16.710 47.960 ;
        RECT 16.980 47.920 17.400 48.200 ;
        RECT 18.620 48.090 18.790 48.420 ;
        RECT 20.240 48.130 20.500 48.220 ;
        RECT 21.150 48.130 21.410 48.220 ;
        RECT 17.920 47.920 19.340 48.090 ;
        RECT 20.150 47.920 20.570 48.130 ;
        RECT 21.080 47.920 21.500 48.130 ;
        RECT 16.980 47.480 18.560 47.650 ;
        RECT 19.770 47.530 19.940 47.860 ;
        RECT 13.810 46.710 13.980 47.040 ;
        RECT 15.220 46.920 16.800 47.090 ;
        RECT 12.280 46.440 12.700 46.650 ;
        RECT 13.170 46.440 13.590 46.650 ;
        RECT 14.400 46.480 15.860 46.650 ;
        RECT 12.350 46.380 12.610 46.440 ;
        RECT 13.260 46.380 13.520 46.440 ;
        RECT 14.860 46.420 15.150 46.480 ;
        RECT 16.380 46.310 16.800 46.650 ;
        RECT 17.060 46.610 17.230 47.480 ;
        RECT 17.610 46.610 17.780 47.300 ;
        RECT 21.750 47.260 21.920 47.950 ;
        RECT 22.290 47.090 22.460 47.960 ;
        RECT 22.730 47.920 23.150 48.200 ;
        RECT 24.370 48.090 24.540 48.420 ;
        RECT 25.990 48.130 26.250 48.220 ;
        RECT 26.900 48.130 27.160 48.220 ;
        RECT 23.670 47.920 25.090 48.090 ;
        RECT 25.900 47.920 26.320 48.130 ;
        RECT 26.830 47.920 27.250 48.130 ;
        RECT 22.730 47.480 24.310 47.650 ;
        RECT 25.520 47.530 25.690 47.860 ;
        RECT 19.560 46.710 19.730 47.040 ;
        RECT 20.970 46.920 22.550 47.090 ;
        RECT 18.030 46.440 18.450 46.650 ;
        RECT 18.920 46.440 19.340 46.650 ;
        RECT 20.150 46.480 21.610 46.650 ;
        RECT 18.100 46.380 18.360 46.440 ;
        RECT 19.010 46.380 19.270 46.440 ;
        RECT 20.610 46.420 20.900 46.480 ;
        RECT 22.130 46.310 22.550 46.650 ;
        RECT 22.810 46.610 22.980 47.480 ;
        RECT 23.360 46.610 23.530 47.300 ;
        RECT 27.500 47.260 27.670 47.950 ;
        RECT 28.040 47.090 28.210 47.960 ;
        RECT 28.480 47.920 28.900 48.200 ;
        RECT 30.120 48.090 30.290 48.420 ;
        RECT 31.740 48.130 32.000 48.220 ;
        RECT 32.650 48.130 32.910 48.220 ;
        RECT 29.420 47.920 30.840 48.090 ;
        RECT 31.650 47.920 32.070 48.130 ;
        RECT 32.580 47.920 33.000 48.130 ;
        RECT 28.480 47.480 30.060 47.650 ;
        RECT 31.270 47.530 31.440 47.860 ;
        RECT 25.310 46.710 25.480 47.040 ;
        RECT 26.720 46.920 28.300 47.090 ;
        RECT 23.780 46.440 24.200 46.650 ;
        RECT 24.670 46.440 25.090 46.650 ;
        RECT 25.900 46.480 27.360 46.650 ;
        RECT 23.850 46.380 24.110 46.440 ;
        RECT 24.760 46.380 25.020 46.440 ;
        RECT 26.360 46.420 26.650 46.480 ;
        RECT 27.880 46.310 28.300 46.650 ;
        RECT 28.560 46.610 28.730 47.480 ;
        RECT 29.110 46.610 29.280 47.300 ;
        RECT 33.250 47.260 33.420 47.950 ;
        RECT 33.790 47.090 33.960 47.960 ;
        RECT 34.230 47.920 34.650 48.200 ;
        RECT 35.870 48.090 36.040 48.420 ;
        RECT 37.490 48.130 37.750 48.220 ;
        RECT 38.400 48.130 38.660 48.220 ;
        RECT 35.170 47.920 36.590 48.090 ;
        RECT 37.400 47.920 37.820 48.130 ;
        RECT 38.330 47.920 38.750 48.130 ;
        RECT 34.230 47.480 35.810 47.650 ;
        RECT 37.020 47.530 37.190 47.860 ;
        RECT 31.060 46.710 31.230 47.040 ;
        RECT 32.470 46.920 34.050 47.090 ;
        RECT 29.530 46.440 29.950 46.650 ;
        RECT 30.420 46.440 30.840 46.650 ;
        RECT 31.650 46.480 33.110 46.650 ;
        RECT 29.600 46.380 29.860 46.440 ;
        RECT 30.510 46.380 30.770 46.440 ;
        RECT 32.110 46.420 32.400 46.480 ;
        RECT 33.630 46.310 34.050 46.650 ;
        RECT 34.310 46.610 34.480 47.480 ;
        RECT 34.860 46.610 35.030 47.300 ;
        RECT 39.000 47.260 39.170 47.950 ;
        RECT 39.540 47.090 39.710 47.960 ;
        RECT 39.980 47.920 40.400 48.200 ;
        RECT 41.620 48.090 41.790 48.420 ;
        RECT 43.240 48.130 43.500 48.220 ;
        RECT 44.150 48.130 44.410 48.220 ;
        RECT 40.920 47.920 42.340 48.090 ;
        RECT 43.150 47.920 43.570 48.130 ;
        RECT 44.080 47.920 44.500 48.130 ;
        RECT 39.980 47.480 41.560 47.650 ;
        RECT 42.770 47.530 42.940 47.860 ;
        RECT 36.810 46.710 36.980 47.040 ;
        RECT 38.220 46.920 39.800 47.090 ;
        RECT 35.280 46.440 35.700 46.650 ;
        RECT 36.170 46.440 36.590 46.650 ;
        RECT 37.400 46.480 38.860 46.650 ;
        RECT 35.350 46.380 35.610 46.440 ;
        RECT 36.260 46.380 36.520 46.440 ;
        RECT 37.860 46.420 38.150 46.480 ;
        RECT 39.380 46.310 39.800 46.650 ;
        RECT 40.060 46.610 40.230 47.480 ;
        RECT 40.610 46.610 40.780 47.300 ;
        RECT 44.750 47.260 44.920 47.950 ;
        RECT 45.290 47.090 45.460 47.960 ;
        RECT 45.730 47.920 46.150 48.200 ;
        RECT 47.370 48.090 47.540 48.420 ;
        RECT 48.990 48.130 49.250 48.220 ;
        RECT 49.900 48.130 50.160 48.220 ;
        RECT 46.670 47.920 48.090 48.090 ;
        RECT 48.900 47.920 49.320 48.130 ;
        RECT 49.830 47.920 50.250 48.130 ;
        RECT 45.730 47.480 47.310 47.650 ;
        RECT 48.520 47.530 48.690 47.860 ;
        RECT 42.560 46.710 42.730 47.040 ;
        RECT 43.970 46.920 45.550 47.090 ;
        RECT 41.030 46.440 41.450 46.650 ;
        RECT 41.920 46.440 42.340 46.650 ;
        RECT 43.150 46.480 44.610 46.650 ;
        RECT 41.100 46.380 41.360 46.440 ;
        RECT 42.010 46.380 42.270 46.440 ;
        RECT 43.610 46.420 43.900 46.480 ;
        RECT 45.130 46.310 45.550 46.650 ;
        RECT 45.810 46.610 45.980 47.480 ;
        RECT 46.360 46.610 46.530 47.300 ;
        RECT 50.500 47.260 50.670 47.950 ;
        RECT 51.040 47.090 51.210 47.960 ;
        RECT 51.480 47.920 51.900 48.200 ;
        RECT 53.120 48.090 53.290 48.420 ;
        RECT 54.740 48.130 55.000 48.220 ;
        RECT 55.650 48.130 55.910 48.220 ;
        RECT 52.420 47.920 53.840 48.090 ;
        RECT 54.650 47.920 55.070 48.130 ;
        RECT 55.580 47.920 56.000 48.130 ;
        RECT 51.480 47.480 53.060 47.650 ;
        RECT 54.270 47.530 54.440 47.860 ;
        RECT 48.310 46.710 48.480 47.040 ;
        RECT 49.720 46.920 51.300 47.090 ;
        RECT 46.780 46.440 47.200 46.650 ;
        RECT 47.670 46.440 48.090 46.650 ;
        RECT 48.900 46.480 50.360 46.650 ;
        RECT 46.850 46.380 47.110 46.440 ;
        RECT 47.760 46.380 48.020 46.440 ;
        RECT 49.360 46.420 49.650 46.480 ;
        RECT 50.880 46.310 51.300 46.650 ;
        RECT 51.560 46.610 51.730 47.480 ;
        RECT 52.110 46.610 52.280 47.300 ;
        RECT 56.250 47.260 56.420 47.950 ;
        RECT 56.790 47.090 56.960 47.960 ;
        RECT 57.230 47.920 57.650 48.200 ;
        RECT 58.870 48.090 59.040 48.420 ;
        RECT 60.490 48.130 60.750 48.220 ;
        RECT 61.400 48.130 61.660 48.220 ;
        RECT 58.170 47.920 59.590 48.090 ;
        RECT 60.400 47.920 60.820 48.130 ;
        RECT 61.330 47.920 61.750 48.130 ;
        RECT 57.230 47.480 58.810 47.650 ;
        RECT 60.020 47.530 60.190 47.860 ;
        RECT 54.060 46.710 54.230 47.040 ;
        RECT 55.470 46.920 57.050 47.090 ;
        RECT 52.530 46.440 52.950 46.650 ;
        RECT 53.420 46.440 53.840 46.650 ;
        RECT 54.650 46.480 56.110 46.650 ;
        RECT 52.600 46.380 52.860 46.440 ;
        RECT 53.510 46.380 53.770 46.440 ;
        RECT 55.110 46.420 55.400 46.480 ;
        RECT 56.630 46.310 57.050 46.650 ;
        RECT 57.310 46.610 57.480 47.480 ;
        RECT 57.860 46.610 58.030 47.300 ;
        RECT 62.000 47.260 62.170 47.950 ;
        RECT 62.540 47.090 62.710 47.960 ;
        RECT 62.980 47.920 63.400 48.200 ;
        RECT 64.620 48.090 64.790 48.420 ;
        RECT 66.240 48.130 66.500 48.220 ;
        RECT 67.150 48.130 67.410 48.220 ;
        RECT 63.920 47.920 65.340 48.090 ;
        RECT 66.150 47.920 66.570 48.130 ;
        RECT 67.080 47.920 67.500 48.130 ;
        RECT 62.980 47.480 64.560 47.650 ;
        RECT 65.770 47.530 65.940 47.860 ;
        RECT 59.810 46.710 59.980 47.040 ;
        RECT 61.220 46.920 62.800 47.090 ;
        RECT 58.280 46.440 58.700 46.650 ;
        RECT 59.170 46.440 59.590 46.650 ;
        RECT 60.400 46.480 61.860 46.650 ;
        RECT 58.350 46.380 58.610 46.440 ;
        RECT 59.260 46.380 59.520 46.440 ;
        RECT 60.860 46.420 61.150 46.480 ;
        RECT 62.380 46.310 62.800 46.650 ;
        RECT 63.060 46.610 63.230 47.480 ;
        RECT 63.610 46.610 63.780 47.300 ;
        RECT 67.750 47.260 67.920 47.950 ;
        RECT 68.290 47.090 68.460 47.960 ;
        RECT 68.730 47.920 69.150 48.200 ;
        RECT 70.370 48.090 70.540 48.420 ;
        RECT 71.990 48.130 72.250 48.220 ;
        RECT 72.900 48.130 73.160 48.220 ;
        RECT 69.670 47.920 71.090 48.090 ;
        RECT 71.900 47.920 72.320 48.130 ;
        RECT 72.830 47.920 73.250 48.130 ;
        RECT 68.730 47.480 70.310 47.650 ;
        RECT 71.520 47.530 71.690 47.860 ;
        RECT 65.560 46.710 65.730 47.040 ;
        RECT 66.970 46.920 68.550 47.090 ;
        RECT 64.030 46.440 64.450 46.650 ;
        RECT 64.920 46.440 65.340 46.650 ;
        RECT 66.150 46.480 67.610 46.650 ;
        RECT 64.100 46.380 64.360 46.440 ;
        RECT 65.010 46.380 65.270 46.440 ;
        RECT 66.610 46.420 66.900 46.480 ;
        RECT 68.130 46.310 68.550 46.650 ;
        RECT 68.810 46.610 68.980 47.480 ;
        RECT 69.360 46.610 69.530 47.300 ;
        RECT 73.500 47.260 73.670 47.950 ;
        RECT 74.040 47.090 74.210 47.960 ;
        RECT 74.480 47.920 74.900 48.200 ;
        RECT 76.120 48.090 76.290 48.420 ;
        RECT 77.740 48.130 78.000 48.220 ;
        RECT 78.650 48.130 78.910 48.220 ;
        RECT 75.420 47.920 76.840 48.090 ;
        RECT 77.650 47.920 78.070 48.130 ;
        RECT 78.580 47.920 79.000 48.130 ;
        RECT 74.480 47.480 76.060 47.650 ;
        RECT 77.270 47.530 77.440 47.860 ;
        RECT 71.310 46.710 71.480 47.040 ;
        RECT 72.720 46.920 74.300 47.090 ;
        RECT 69.780 46.440 70.200 46.650 ;
        RECT 70.670 46.440 71.090 46.650 ;
        RECT 71.900 46.480 73.360 46.650 ;
        RECT 69.850 46.380 70.110 46.440 ;
        RECT 70.760 46.380 71.020 46.440 ;
        RECT 72.360 46.420 72.650 46.480 ;
        RECT 73.880 46.310 74.300 46.650 ;
        RECT 74.560 46.610 74.730 47.480 ;
        RECT 75.110 46.610 75.280 47.300 ;
        RECT 79.250 47.260 79.420 47.950 ;
        RECT 79.790 47.090 79.960 47.960 ;
        RECT 80.230 47.920 80.650 48.200 ;
        RECT 81.870 48.090 82.040 48.420 ;
        RECT 83.490 48.130 83.750 48.220 ;
        RECT 84.400 48.130 84.660 48.220 ;
        RECT 81.170 47.920 82.590 48.090 ;
        RECT 83.400 47.920 83.820 48.130 ;
        RECT 84.330 47.920 84.750 48.130 ;
        RECT 80.230 47.480 81.810 47.650 ;
        RECT 83.020 47.530 83.190 47.860 ;
        RECT 77.060 46.710 77.230 47.040 ;
        RECT 78.470 46.920 80.050 47.090 ;
        RECT 75.530 46.440 75.950 46.650 ;
        RECT 76.420 46.440 76.840 46.650 ;
        RECT 77.650 46.480 79.110 46.650 ;
        RECT 75.600 46.380 75.860 46.440 ;
        RECT 76.510 46.380 76.770 46.440 ;
        RECT 78.110 46.420 78.400 46.480 ;
        RECT 79.630 46.310 80.050 46.650 ;
        RECT 80.310 46.610 80.480 47.480 ;
        RECT 80.860 46.610 81.030 47.300 ;
        RECT 85.000 47.260 85.170 47.950 ;
        RECT 85.540 47.090 85.710 47.960 ;
        RECT 85.980 47.920 86.400 48.200 ;
        RECT 87.620 48.090 87.790 48.420 ;
        RECT 89.240 48.130 89.500 48.220 ;
        RECT 90.150 48.130 90.410 48.220 ;
        RECT 86.920 47.920 88.340 48.090 ;
        RECT 89.150 47.920 89.570 48.130 ;
        RECT 90.080 47.920 90.500 48.130 ;
        RECT 85.980 47.480 87.560 47.650 ;
        RECT 88.770 47.530 88.940 47.860 ;
        RECT 82.810 46.710 82.980 47.040 ;
        RECT 84.220 46.920 85.800 47.090 ;
        RECT 81.280 46.440 81.700 46.650 ;
        RECT 82.170 46.440 82.590 46.650 ;
        RECT 83.400 46.480 84.860 46.650 ;
        RECT 81.350 46.380 81.610 46.440 ;
        RECT 82.260 46.380 82.520 46.440 ;
        RECT 83.860 46.420 84.150 46.480 ;
        RECT 85.380 46.310 85.800 46.650 ;
        RECT 86.060 46.610 86.230 47.480 ;
        RECT 86.610 46.610 86.780 47.300 ;
        RECT 90.750 47.260 90.920 47.950 ;
        RECT 91.290 47.090 91.460 47.960 ;
        RECT 91.730 47.920 92.150 48.200 ;
        RECT 93.370 48.090 93.540 48.420 ;
        RECT 92.670 47.920 94.090 48.090 ;
        RECT 91.730 47.480 93.310 47.650 ;
        RECT 88.560 46.710 88.730 47.040 ;
        RECT 89.970 46.920 91.550 47.090 ;
        RECT 87.030 46.440 87.450 46.650 ;
        RECT 87.920 46.440 88.340 46.650 ;
        RECT 89.150 46.480 90.610 46.650 ;
        RECT 87.100 46.380 87.360 46.440 ;
        RECT 88.010 46.380 88.270 46.440 ;
        RECT 89.610 46.420 89.900 46.480 ;
        RECT 91.130 46.310 91.550 46.650 ;
        RECT 91.810 46.610 91.980 47.480 ;
        RECT 92.360 46.610 92.530 47.300 ;
        RECT 94.310 46.710 94.480 47.040 ;
        RECT 92.780 46.440 93.200 46.650 ;
        RECT 93.670 46.440 94.090 46.650 ;
        RECT 92.850 46.380 93.110 46.440 ;
        RECT 93.760 46.380 94.020 46.440 ;
        RECT 2.990 45.720 3.250 45.810 ;
        RECT 3.900 45.720 4.160 45.810 ;
        RECT 2.900 45.510 3.320 45.720 ;
        RECT 3.830 45.510 4.250 45.720 ;
        RECT 2.520 45.120 2.690 45.450 ;
        RECT 4.500 44.850 4.670 45.540 ;
        RECT 5.040 44.680 5.210 45.550 ;
        RECT 5.480 45.510 5.900 45.790 ;
        RECT 7.120 45.680 7.290 46.010 ;
        RECT 8.740 45.720 9.000 45.810 ;
        RECT 9.650 45.720 9.910 45.810 ;
        RECT 6.420 45.510 7.840 45.680 ;
        RECT 8.650 45.510 9.070 45.720 ;
        RECT 9.580 45.510 10.000 45.720 ;
        RECT 5.480 45.070 7.060 45.240 ;
        RECT 8.270 45.120 8.440 45.450 ;
        RECT 3.720 44.510 5.300 44.680 ;
        RECT 2.900 44.070 4.360 44.240 ;
        RECT 3.020 43.190 3.190 44.070 ;
        RECT 3.360 44.010 3.650 44.070 ;
        RECT 4.880 43.900 5.300 44.240 ;
        RECT 5.560 44.200 5.730 45.070 ;
        RECT 6.110 44.200 6.280 44.890 ;
        RECT 10.250 44.850 10.420 45.540 ;
        RECT 10.790 44.680 10.960 45.550 ;
        RECT 11.230 45.510 11.650 45.790 ;
        RECT 12.870 45.680 13.040 46.010 ;
        RECT 14.490 45.720 14.750 45.810 ;
        RECT 15.400 45.720 15.660 45.810 ;
        RECT 12.170 45.510 13.590 45.680 ;
        RECT 14.400 45.510 14.820 45.720 ;
        RECT 15.330 45.510 15.750 45.720 ;
        RECT 11.230 45.070 12.810 45.240 ;
        RECT 14.020 45.120 14.190 45.450 ;
        RECT 8.060 44.300 8.230 44.630 ;
        RECT 9.470 44.510 11.050 44.680 ;
        RECT 6.530 44.030 6.950 44.240 ;
        RECT 7.420 44.030 7.840 44.240 ;
        RECT 8.650 44.070 10.110 44.240 ;
        RECT 6.600 43.970 6.860 44.030 ;
        RECT 7.510 43.970 7.770 44.030 ;
        RECT 5.010 43.190 5.180 43.900 ;
        RECT 2.990 42.750 3.250 42.840 ;
        RECT 3.900 42.750 4.160 42.840 ;
        RECT 2.900 42.540 3.320 42.750 ;
        RECT 3.830 42.540 4.250 42.750 ;
        RECT 2.520 42.150 2.690 42.480 ;
        RECT 4.500 41.880 4.670 42.570 ;
        RECT 5.040 41.710 5.210 42.580 ;
        RECT 5.480 42.540 5.900 42.820 ;
        RECT 7.120 42.710 7.290 43.280 ;
        RECT 8.770 43.190 8.940 44.070 ;
        RECT 9.110 44.010 9.400 44.070 ;
        RECT 10.630 43.900 11.050 44.240 ;
        RECT 11.310 44.200 11.480 45.070 ;
        RECT 11.860 44.200 12.030 44.890 ;
        RECT 16.000 44.850 16.170 45.540 ;
        RECT 16.540 44.680 16.710 45.550 ;
        RECT 16.980 45.510 17.400 45.790 ;
        RECT 18.620 45.680 18.790 46.010 ;
        RECT 20.240 45.720 20.500 45.810 ;
        RECT 21.150 45.720 21.410 45.810 ;
        RECT 17.920 45.510 19.340 45.680 ;
        RECT 20.150 45.510 20.570 45.720 ;
        RECT 21.080 45.510 21.500 45.720 ;
        RECT 16.980 45.070 18.560 45.240 ;
        RECT 19.770 45.120 19.940 45.450 ;
        RECT 13.810 44.300 13.980 44.630 ;
        RECT 15.220 44.510 16.800 44.680 ;
        RECT 12.280 44.030 12.700 44.240 ;
        RECT 13.170 44.030 13.590 44.240 ;
        RECT 14.400 44.070 15.860 44.240 ;
        RECT 12.350 43.970 12.610 44.030 ;
        RECT 13.260 43.970 13.520 44.030 ;
        RECT 10.770 43.190 10.940 43.900 ;
        RECT 8.740 42.750 9.000 42.840 ;
        RECT 9.650 42.750 9.910 42.840 ;
        RECT 6.420 42.540 7.840 42.710 ;
        RECT 8.650 42.540 9.070 42.750 ;
        RECT 9.580 42.540 10.000 42.750 ;
        RECT 5.480 42.100 7.060 42.270 ;
        RECT 8.270 42.150 8.440 42.480 ;
        RECT 3.720 41.540 5.300 41.710 ;
        RECT 2.900 41.100 4.360 41.270 ;
        RECT 3.360 41.040 3.650 41.100 ;
        RECT 4.880 40.930 5.300 41.270 ;
        RECT 5.560 41.230 5.730 42.100 ;
        RECT 6.110 41.230 6.280 41.920 ;
        RECT 10.250 41.880 10.420 42.570 ;
        RECT 10.790 41.710 10.960 42.580 ;
        RECT 11.230 42.540 11.650 42.820 ;
        RECT 12.870 42.710 13.040 43.280 ;
        RECT 14.520 43.190 14.690 44.070 ;
        RECT 14.860 44.010 15.150 44.070 ;
        RECT 16.380 43.900 16.800 44.240 ;
        RECT 17.060 44.200 17.230 45.070 ;
        RECT 17.610 44.200 17.780 44.890 ;
        RECT 21.750 44.850 21.920 45.540 ;
        RECT 22.290 44.680 22.460 45.550 ;
        RECT 22.730 45.510 23.150 45.790 ;
        RECT 24.370 45.680 24.540 46.010 ;
        RECT 25.990 45.720 26.250 45.810 ;
        RECT 26.900 45.720 27.160 45.810 ;
        RECT 23.670 45.510 25.090 45.680 ;
        RECT 25.900 45.510 26.320 45.720 ;
        RECT 26.830 45.510 27.250 45.720 ;
        RECT 22.730 45.070 24.310 45.240 ;
        RECT 25.520 45.120 25.690 45.450 ;
        RECT 19.560 44.300 19.730 44.630 ;
        RECT 20.970 44.510 22.550 44.680 ;
        RECT 18.030 44.030 18.450 44.240 ;
        RECT 18.920 44.030 19.340 44.240 ;
        RECT 20.150 44.070 21.610 44.240 ;
        RECT 18.100 43.970 18.360 44.030 ;
        RECT 19.010 43.970 19.270 44.030 ;
        RECT 16.520 43.190 16.690 43.900 ;
        RECT 14.490 42.750 14.750 42.840 ;
        RECT 15.400 42.750 15.660 42.840 ;
        RECT 12.170 42.540 13.590 42.710 ;
        RECT 14.400 42.540 14.820 42.750 ;
        RECT 15.330 42.540 15.750 42.750 ;
        RECT 11.230 42.100 12.810 42.270 ;
        RECT 14.020 42.150 14.190 42.480 ;
        RECT 8.060 41.330 8.230 41.660 ;
        RECT 9.470 41.540 11.050 41.710 ;
        RECT 6.530 41.060 6.950 41.270 ;
        RECT 7.420 41.060 7.840 41.270 ;
        RECT 8.650 41.100 10.110 41.270 ;
        RECT 6.600 41.000 6.860 41.060 ;
        RECT 7.510 41.000 7.770 41.060 ;
        RECT 9.110 41.040 9.400 41.100 ;
        RECT 10.630 40.930 11.050 41.270 ;
        RECT 11.310 41.230 11.480 42.100 ;
        RECT 11.860 41.230 12.030 41.920 ;
        RECT 16.000 41.880 16.170 42.570 ;
        RECT 16.540 41.710 16.710 42.580 ;
        RECT 16.980 42.540 17.400 42.820 ;
        RECT 18.620 42.710 18.790 43.280 ;
        RECT 20.270 43.190 20.440 44.070 ;
        RECT 20.610 44.010 20.900 44.070 ;
        RECT 22.130 43.900 22.550 44.240 ;
        RECT 22.810 44.200 22.980 45.070 ;
        RECT 23.360 44.200 23.530 44.890 ;
        RECT 27.500 44.850 27.670 45.540 ;
        RECT 28.040 44.680 28.210 45.550 ;
        RECT 28.480 45.510 28.900 45.790 ;
        RECT 30.120 45.680 30.290 46.010 ;
        RECT 31.740 45.720 32.000 45.810 ;
        RECT 32.650 45.720 32.910 45.810 ;
        RECT 29.420 45.510 30.840 45.680 ;
        RECT 31.650 45.510 32.070 45.720 ;
        RECT 32.580 45.510 33.000 45.720 ;
        RECT 28.480 45.070 30.060 45.240 ;
        RECT 31.270 45.120 31.440 45.450 ;
        RECT 25.310 44.300 25.480 44.630 ;
        RECT 26.720 44.510 28.300 44.680 ;
        RECT 23.780 44.030 24.200 44.240 ;
        RECT 24.670 44.030 25.090 44.240 ;
        RECT 25.900 44.070 27.360 44.240 ;
        RECT 23.850 43.970 24.110 44.030 ;
        RECT 24.760 43.970 25.020 44.030 ;
        RECT 22.270 43.190 22.440 43.900 ;
        RECT 20.240 42.750 20.500 42.840 ;
        RECT 21.150 42.750 21.410 42.840 ;
        RECT 17.920 42.540 19.340 42.710 ;
        RECT 20.150 42.540 20.570 42.750 ;
        RECT 21.080 42.540 21.500 42.750 ;
        RECT 16.980 42.100 18.560 42.270 ;
        RECT 19.770 42.150 19.940 42.480 ;
        RECT 13.810 41.330 13.980 41.660 ;
        RECT 15.220 41.540 16.800 41.710 ;
        RECT 12.280 41.060 12.700 41.270 ;
        RECT 13.170 41.060 13.590 41.270 ;
        RECT 14.400 41.100 15.860 41.270 ;
        RECT 12.350 41.000 12.610 41.060 ;
        RECT 13.260 41.000 13.520 41.060 ;
        RECT 14.860 41.040 15.150 41.100 ;
        RECT 16.380 40.930 16.800 41.270 ;
        RECT 17.060 41.230 17.230 42.100 ;
        RECT 17.610 41.230 17.780 41.920 ;
        RECT 21.750 41.880 21.920 42.570 ;
        RECT 22.290 41.710 22.460 42.580 ;
        RECT 22.730 42.540 23.150 42.820 ;
        RECT 24.370 42.710 24.540 43.280 ;
        RECT 26.020 43.190 26.190 44.070 ;
        RECT 26.360 44.010 26.650 44.070 ;
        RECT 27.880 43.900 28.300 44.240 ;
        RECT 28.560 44.200 28.730 45.070 ;
        RECT 29.110 44.200 29.280 44.890 ;
        RECT 33.250 44.850 33.420 45.540 ;
        RECT 33.790 44.680 33.960 45.550 ;
        RECT 34.230 45.510 34.650 45.790 ;
        RECT 35.870 45.680 36.040 46.010 ;
        RECT 37.490 45.720 37.750 45.810 ;
        RECT 38.400 45.720 38.660 45.810 ;
        RECT 35.170 45.510 36.590 45.680 ;
        RECT 37.400 45.510 37.820 45.720 ;
        RECT 38.330 45.510 38.750 45.720 ;
        RECT 34.230 45.070 35.810 45.240 ;
        RECT 37.020 45.120 37.190 45.450 ;
        RECT 31.060 44.300 31.230 44.630 ;
        RECT 32.470 44.510 34.050 44.680 ;
        RECT 29.530 44.030 29.950 44.240 ;
        RECT 30.420 44.030 30.840 44.240 ;
        RECT 31.650 44.070 33.110 44.240 ;
        RECT 29.600 43.970 29.860 44.030 ;
        RECT 30.510 43.970 30.770 44.030 ;
        RECT 28.020 43.190 28.190 43.900 ;
        RECT 25.990 42.750 26.250 42.840 ;
        RECT 26.900 42.750 27.160 42.840 ;
        RECT 23.670 42.540 25.090 42.710 ;
        RECT 25.900 42.540 26.320 42.750 ;
        RECT 26.830 42.540 27.250 42.750 ;
        RECT 22.730 42.100 24.310 42.270 ;
        RECT 25.520 42.150 25.690 42.480 ;
        RECT 19.560 41.330 19.730 41.660 ;
        RECT 20.970 41.540 22.550 41.710 ;
        RECT 18.030 41.060 18.450 41.270 ;
        RECT 18.920 41.060 19.340 41.270 ;
        RECT 20.150 41.100 21.610 41.270 ;
        RECT 18.100 41.000 18.360 41.060 ;
        RECT 19.010 41.000 19.270 41.060 ;
        RECT 20.610 41.040 20.900 41.100 ;
        RECT 22.130 40.930 22.550 41.270 ;
        RECT 22.810 41.230 22.980 42.100 ;
        RECT 23.360 41.230 23.530 41.920 ;
        RECT 27.500 41.880 27.670 42.570 ;
        RECT 28.040 41.710 28.210 42.580 ;
        RECT 28.480 42.540 28.900 42.820 ;
        RECT 30.120 42.710 30.290 43.280 ;
        RECT 31.770 43.190 31.940 44.070 ;
        RECT 32.110 44.010 32.400 44.070 ;
        RECT 33.630 43.900 34.050 44.240 ;
        RECT 34.310 44.200 34.480 45.070 ;
        RECT 34.860 44.200 35.030 44.890 ;
        RECT 39.000 44.850 39.170 45.540 ;
        RECT 39.540 44.680 39.710 45.550 ;
        RECT 39.980 45.510 40.400 45.790 ;
        RECT 41.620 45.680 41.790 46.010 ;
        RECT 43.240 45.720 43.500 45.810 ;
        RECT 44.150 45.720 44.410 45.810 ;
        RECT 40.920 45.510 42.340 45.680 ;
        RECT 43.150 45.510 43.570 45.720 ;
        RECT 44.080 45.510 44.500 45.720 ;
        RECT 39.980 45.070 41.560 45.240 ;
        RECT 42.770 45.120 42.940 45.450 ;
        RECT 36.810 44.300 36.980 44.630 ;
        RECT 38.220 44.510 39.800 44.680 ;
        RECT 35.280 44.030 35.700 44.240 ;
        RECT 36.170 44.030 36.590 44.240 ;
        RECT 37.400 44.070 38.860 44.240 ;
        RECT 35.350 43.970 35.610 44.030 ;
        RECT 36.260 43.970 36.520 44.030 ;
        RECT 33.770 43.190 33.940 43.900 ;
        RECT 31.740 42.750 32.000 42.840 ;
        RECT 32.650 42.750 32.910 42.840 ;
        RECT 29.420 42.540 30.840 42.710 ;
        RECT 31.650 42.540 32.070 42.750 ;
        RECT 32.580 42.540 33.000 42.750 ;
        RECT 28.480 42.100 30.060 42.270 ;
        RECT 31.270 42.150 31.440 42.480 ;
        RECT 25.310 41.330 25.480 41.660 ;
        RECT 26.720 41.540 28.300 41.710 ;
        RECT 23.780 41.060 24.200 41.270 ;
        RECT 24.670 41.060 25.090 41.270 ;
        RECT 25.900 41.100 27.360 41.270 ;
        RECT 23.850 41.000 24.110 41.060 ;
        RECT 24.760 41.000 25.020 41.060 ;
        RECT 26.360 41.040 26.650 41.100 ;
        RECT 27.880 40.930 28.300 41.270 ;
        RECT 28.560 41.230 28.730 42.100 ;
        RECT 29.110 41.230 29.280 41.920 ;
        RECT 33.250 41.880 33.420 42.570 ;
        RECT 33.790 41.710 33.960 42.580 ;
        RECT 34.230 42.540 34.650 42.820 ;
        RECT 35.870 42.710 36.040 43.280 ;
        RECT 37.520 43.190 37.690 44.070 ;
        RECT 37.860 44.010 38.150 44.070 ;
        RECT 39.380 43.900 39.800 44.240 ;
        RECT 40.060 44.200 40.230 45.070 ;
        RECT 40.610 44.200 40.780 44.890 ;
        RECT 44.750 44.850 44.920 45.540 ;
        RECT 45.290 44.680 45.460 45.550 ;
        RECT 45.730 45.510 46.150 45.790 ;
        RECT 47.370 45.680 47.540 46.010 ;
        RECT 48.990 45.720 49.250 45.810 ;
        RECT 49.900 45.720 50.160 45.810 ;
        RECT 46.670 45.510 48.090 45.680 ;
        RECT 48.900 45.510 49.320 45.720 ;
        RECT 49.830 45.510 50.250 45.720 ;
        RECT 45.730 45.070 47.310 45.240 ;
        RECT 48.520 45.120 48.690 45.450 ;
        RECT 42.560 44.300 42.730 44.630 ;
        RECT 43.970 44.510 45.550 44.680 ;
        RECT 41.030 44.030 41.450 44.240 ;
        RECT 41.920 44.030 42.340 44.240 ;
        RECT 43.150 44.070 44.610 44.240 ;
        RECT 41.100 43.970 41.360 44.030 ;
        RECT 42.010 43.970 42.270 44.030 ;
        RECT 39.520 43.190 39.690 43.900 ;
        RECT 37.490 42.750 37.750 42.840 ;
        RECT 38.400 42.750 38.660 42.840 ;
        RECT 35.170 42.540 36.590 42.710 ;
        RECT 37.400 42.540 37.820 42.750 ;
        RECT 38.330 42.540 38.750 42.750 ;
        RECT 34.230 42.100 35.810 42.270 ;
        RECT 37.020 42.150 37.190 42.480 ;
        RECT 31.060 41.330 31.230 41.660 ;
        RECT 32.470 41.540 34.050 41.710 ;
        RECT 29.530 41.060 29.950 41.270 ;
        RECT 30.420 41.060 30.840 41.270 ;
        RECT 31.650 41.100 33.110 41.270 ;
        RECT 29.600 41.000 29.860 41.060 ;
        RECT 30.510 41.000 30.770 41.060 ;
        RECT 32.110 41.040 32.400 41.100 ;
        RECT 33.630 40.930 34.050 41.270 ;
        RECT 34.310 41.230 34.480 42.100 ;
        RECT 34.860 41.230 35.030 41.920 ;
        RECT 39.000 41.880 39.170 42.570 ;
        RECT 39.540 41.710 39.710 42.580 ;
        RECT 39.980 42.540 40.400 42.820 ;
        RECT 41.620 42.710 41.790 43.280 ;
        RECT 43.270 43.190 43.440 44.070 ;
        RECT 43.610 44.010 43.900 44.070 ;
        RECT 45.130 43.900 45.550 44.240 ;
        RECT 45.810 44.200 45.980 45.070 ;
        RECT 46.360 44.200 46.530 44.890 ;
        RECT 50.500 44.850 50.670 45.540 ;
        RECT 51.040 44.680 51.210 45.550 ;
        RECT 51.480 45.510 51.900 45.790 ;
        RECT 53.120 45.680 53.290 46.010 ;
        RECT 54.740 45.720 55.000 45.810 ;
        RECT 55.650 45.720 55.910 45.810 ;
        RECT 52.420 45.510 53.840 45.680 ;
        RECT 54.650 45.510 55.070 45.720 ;
        RECT 55.580 45.510 56.000 45.720 ;
        RECT 51.480 45.070 53.060 45.240 ;
        RECT 54.270 45.120 54.440 45.450 ;
        RECT 48.310 44.300 48.480 44.630 ;
        RECT 49.720 44.510 51.300 44.680 ;
        RECT 46.780 44.030 47.200 44.240 ;
        RECT 47.670 44.030 48.090 44.240 ;
        RECT 48.900 44.070 50.360 44.240 ;
        RECT 46.850 43.970 47.110 44.030 ;
        RECT 47.760 43.970 48.020 44.030 ;
        RECT 45.270 43.190 45.440 43.900 ;
        RECT 43.240 42.750 43.500 42.840 ;
        RECT 44.150 42.750 44.410 42.840 ;
        RECT 40.920 42.540 42.340 42.710 ;
        RECT 43.150 42.540 43.570 42.750 ;
        RECT 44.080 42.540 44.500 42.750 ;
        RECT 39.980 42.100 41.560 42.270 ;
        RECT 42.770 42.150 42.940 42.480 ;
        RECT 36.810 41.330 36.980 41.660 ;
        RECT 38.220 41.540 39.800 41.710 ;
        RECT 35.280 41.060 35.700 41.270 ;
        RECT 36.170 41.060 36.590 41.270 ;
        RECT 37.400 41.100 38.860 41.270 ;
        RECT 35.350 41.000 35.610 41.060 ;
        RECT 36.260 41.000 36.520 41.060 ;
        RECT 37.860 41.040 38.150 41.100 ;
        RECT 39.380 40.930 39.800 41.270 ;
        RECT 40.060 41.230 40.230 42.100 ;
        RECT 40.610 41.230 40.780 41.920 ;
        RECT 44.750 41.880 44.920 42.570 ;
        RECT 45.290 41.710 45.460 42.580 ;
        RECT 45.730 42.540 46.150 42.820 ;
        RECT 47.370 42.710 47.540 43.280 ;
        RECT 49.020 43.190 49.190 44.070 ;
        RECT 49.360 44.010 49.650 44.070 ;
        RECT 50.880 43.900 51.300 44.240 ;
        RECT 51.560 44.200 51.730 45.070 ;
        RECT 52.110 44.200 52.280 44.890 ;
        RECT 56.250 44.850 56.420 45.540 ;
        RECT 56.790 44.680 56.960 45.550 ;
        RECT 57.230 45.510 57.650 45.790 ;
        RECT 58.870 45.680 59.040 46.010 ;
        RECT 60.490 45.720 60.750 45.810 ;
        RECT 61.400 45.720 61.660 45.810 ;
        RECT 58.170 45.510 59.590 45.680 ;
        RECT 60.400 45.510 60.820 45.720 ;
        RECT 61.330 45.510 61.750 45.720 ;
        RECT 57.230 45.070 58.810 45.240 ;
        RECT 60.020 45.120 60.190 45.450 ;
        RECT 54.060 44.300 54.230 44.630 ;
        RECT 55.470 44.510 57.050 44.680 ;
        RECT 52.530 44.030 52.950 44.240 ;
        RECT 53.420 44.030 53.840 44.240 ;
        RECT 54.650 44.070 56.110 44.240 ;
        RECT 52.600 43.970 52.860 44.030 ;
        RECT 53.510 43.970 53.770 44.030 ;
        RECT 51.020 43.190 51.190 43.900 ;
        RECT 48.990 42.750 49.250 42.840 ;
        RECT 49.900 42.750 50.160 42.840 ;
        RECT 46.670 42.540 48.090 42.710 ;
        RECT 48.900 42.540 49.320 42.750 ;
        RECT 49.830 42.540 50.250 42.750 ;
        RECT 45.730 42.100 47.310 42.270 ;
        RECT 48.520 42.150 48.690 42.480 ;
        RECT 42.560 41.330 42.730 41.660 ;
        RECT 43.970 41.540 45.550 41.710 ;
        RECT 41.030 41.060 41.450 41.270 ;
        RECT 41.920 41.060 42.340 41.270 ;
        RECT 43.150 41.100 44.610 41.270 ;
        RECT 41.100 41.000 41.360 41.060 ;
        RECT 42.010 41.000 42.270 41.060 ;
        RECT 43.610 41.040 43.900 41.100 ;
        RECT 45.130 40.930 45.550 41.270 ;
        RECT 45.810 41.230 45.980 42.100 ;
        RECT 46.360 41.230 46.530 41.920 ;
        RECT 50.500 41.880 50.670 42.570 ;
        RECT 51.040 41.710 51.210 42.580 ;
        RECT 51.480 42.540 51.900 42.820 ;
        RECT 53.120 42.710 53.290 43.280 ;
        RECT 54.770 43.190 54.940 44.070 ;
        RECT 55.110 44.010 55.400 44.070 ;
        RECT 56.630 43.900 57.050 44.240 ;
        RECT 57.310 44.200 57.480 45.070 ;
        RECT 57.860 44.200 58.030 44.890 ;
        RECT 62.000 44.850 62.170 45.540 ;
        RECT 62.540 44.680 62.710 45.550 ;
        RECT 62.980 45.510 63.400 45.790 ;
        RECT 64.620 45.680 64.790 46.010 ;
        RECT 66.240 45.720 66.500 45.810 ;
        RECT 67.150 45.720 67.410 45.810 ;
        RECT 63.920 45.510 65.340 45.680 ;
        RECT 66.150 45.510 66.570 45.720 ;
        RECT 67.080 45.510 67.500 45.720 ;
        RECT 62.980 45.070 64.560 45.240 ;
        RECT 65.770 45.120 65.940 45.450 ;
        RECT 59.810 44.300 59.980 44.630 ;
        RECT 61.220 44.510 62.800 44.680 ;
        RECT 58.280 44.030 58.700 44.240 ;
        RECT 59.170 44.030 59.590 44.240 ;
        RECT 60.400 44.070 61.860 44.240 ;
        RECT 58.350 43.970 58.610 44.030 ;
        RECT 59.260 43.970 59.520 44.030 ;
        RECT 56.770 43.190 56.940 43.900 ;
        RECT 54.740 42.750 55.000 42.840 ;
        RECT 55.650 42.750 55.910 42.840 ;
        RECT 52.420 42.540 53.840 42.710 ;
        RECT 54.650 42.540 55.070 42.750 ;
        RECT 55.580 42.540 56.000 42.750 ;
        RECT 51.480 42.100 53.060 42.270 ;
        RECT 54.270 42.150 54.440 42.480 ;
        RECT 48.310 41.330 48.480 41.660 ;
        RECT 49.720 41.540 51.300 41.710 ;
        RECT 46.780 41.060 47.200 41.270 ;
        RECT 47.670 41.060 48.090 41.270 ;
        RECT 48.900 41.100 50.360 41.270 ;
        RECT 46.850 41.000 47.110 41.060 ;
        RECT 47.760 41.000 48.020 41.060 ;
        RECT 49.360 41.040 49.650 41.100 ;
        RECT 50.880 40.930 51.300 41.270 ;
        RECT 51.560 41.230 51.730 42.100 ;
        RECT 52.110 41.230 52.280 41.920 ;
        RECT 56.250 41.880 56.420 42.570 ;
        RECT 56.790 41.710 56.960 42.580 ;
        RECT 57.230 42.540 57.650 42.820 ;
        RECT 58.870 42.710 59.040 43.280 ;
        RECT 60.520 43.190 60.690 44.070 ;
        RECT 60.860 44.010 61.150 44.070 ;
        RECT 62.380 43.900 62.800 44.240 ;
        RECT 63.060 44.200 63.230 45.070 ;
        RECT 63.610 44.200 63.780 44.890 ;
        RECT 67.750 44.850 67.920 45.540 ;
        RECT 68.290 44.680 68.460 45.550 ;
        RECT 68.730 45.510 69.150 45.790 ;
        RECT 70.370 45.680 70.540 46.010 ;
        RECT 71.990 45.720 72.250 45.810 ;
        RECT 72.900 45.720 73.160 45.810 ;
        RECT 69.670 45.510 71.090 45.680 ;
        RECT 71.900 45.510 72.320 45.720 ;
        RECT 72.830 45.510 73.250 45.720 ;
        RECT 68.730 45.070 70.310 45.240 ;
        RECT 71.520 45.120 71.690 45.450 ;
        RECT 65.560 44.300 65.730 44.630 ;
        RECT 66.970 44.510 68.550 44.680 ;
        RECT 64.030 44.030 64.450 44.240 ;
        RECT 64.920 44.030 65.340 44.240 ;
        RECT 66.150 44.070 67.610 44.240 ;
        RECT 64.100 43.970 64.360 44.030 ;
        RECT 65.010 43.970 65.270 44.030 ;
        RECT 62.520 43.190 62.690 43.900 ;
        RECT 60.490 42.750 60.750 42.840 ;
        RECT 61.400 42.750 61.660 42.840 ;
        RECT 58.170 42.540 59.590 42.710 ;
        RECT 60.400 42.540 60.820 42.750 ;
        RECT 61.330 42.540 61.750 42.750 ;
        RECT 57.230 42.100 58.810 42.270 ;
        RECT 60.020 42.150 60.190 42.480 ;
        RECT 54.060 41.330 54.230 41.660 ;
        RECT 55.470 41.540 57.050 41.710 ;
        RECT 52.530 41.060 52.950 41.270 ;
        RECT 53.420 41.060 53.840 41.270 ;
        RECT 54.650 41.100 56.110 41.270 ;
        RECT 52.600 41.000 52.860 41.060 ;
        RECT 53.510 41.000 53.770 41.060 ;
        RECT 55.110 41.040 55.400 41.100 ;
        RECT 56.630 40.930 57.050 41.270 ;
        RECT 57.310 41.230 57.480 42.100 ;
        RECT 57.860 41.230 58.030 41.920 ;
        RECT 62.000 41.880 62.170 42.570 ;
        RECT 62.540 41.710 62.710 42.580 ;
        RECT 62.980 42.540 63.400 42.820 ;
        RECT 64.620 42.710 64.790 43.280 ;
        RECT 66.270 43.190 66.440 44.070 ;
        RECT 66.610 44.010 66.900 44.070 ;
        RECT 68.130 43.900 68.550 44.240 ;
        RECT 68.810 44.200 68.980 45.070 ;
        RECT 69.360 44.200 69.530 44.890 ;
        RECT 73.500 44.850 73.670 45.540 ;
        RECT 74.040 44.680 74.210 45.550 ;
        RECT 74.480 45.510 74.900 45.790 ;
        RECT 76.120 45.680 76.290 46.010 ;
        RECT 77.740 45.720 78.000 45.810 ;
        RECT 78.650 45.720 78.910 45.810 ;
        RECT 75.420 45.510 76.840 45.680 ;
        RECT 77.650 45.510 78.070 45.720 ;
        RECT 78.580 45.510 79.000 45.720 ;
        RECT 74.480 45.070 76.060 45.240 ;
        RECT 77.270 45.120 77.440 45.450 ;
        RECT 71.310 44.300 71.480 44.630 ;
        RECT 72.720 44.510 74.300 44.680 ;
        RECT 69.780 44.030 70.200 44.240 ;
        RECT 70.670 44.030 71.090 44.240 ;
        RECT 71.900 44.070 73.360 44.240 ;
        RECT 69.850 43.970 70.110 44.030 ;
        RECT 70.760 43.970 71.020 44.030 ;
        RECT 68.270 43.190 68.440 43.900 ;
        RECT 66.240 42.750 66.500 42.840 ;
        RECT 67.150 42.750 67.410 42.840 ;
        RECT 63.920 42.540 65.340 42.710 ;
        RECT 66.150 42.540 66.570 42.750 ;
        RECT 67.080 42.540 67.500 42.750 ;
        RECT 62.980 42.100 64.560 42.270 ;
        RECT 65.770 42.150 65.940 42.480 ;
        RECT 59.810 41.330 59.980 41.660 ;
        RECT 61.220 41.540 62.800 41.710 ;
        RECT 58.280 41.060 58.700 41.270 ;
        RECT 59.170 41.060 59.590 41.270 ;
        RECT 60.400 41.100 61.860 41.270 ;
        RECT 58.350 41.000 58.610 41.060 ;
        RECT 59.260 41.000 59.520 41.060 ;
        RECT 60.860 41.040 61.150 41.100 ;
        RECT 62.380 40.930 62.800 41.270 ;
        RECT 63.060 41.230 63.230 42.100 ;
        RECT 63.610 41.230 63.780 41.920 ;
        RECT 67.750 41.880 67.920 42.570 ;
        RECT 68.290 41.710 68.460 42.580 ;
        RECT 68.730 42.540 69.150 42.820 ;
        RECT 70.370 42.710 70.540 43.280 ;
        RECT 72.020 43.190 72.190 44.070 ;
        RECT 72.360 44.010 72.650 44.070 ;
        RECT 73.880 43.900 74.300 44.240 ;
        RECT 74.560 44.200 74.730 45.070 ;
        RECT 75.110 44.200 75.280 44.890 ;
        RECT 79.250 44.850 79.420 45.540 ;
        RECT 79.790 44.680 79.960 45.550 ;
        RECT 80.230 45.510 80.650 45.790 ;
        RECT 81.870 45.680 82.040 46.010 ;
        RECT 83.490 45.720 83.750 45.810 ;
        RECT 84.400 45.720 84.660 45.810 ;
        RECT 81.170 45.510 82.590 45.680 ;
        RECT 83.400 45.510 83.820 45.720 ;
        RECT 84.330 45.510 84.750 45.720 ;
        RECT 80.230 45.070 81.810 45.240 ;
        RECT 83.020 45.120 83.190 45.450 ;
        RECT 77.060 44.300 77.230 44.630 ;
        RECT 78.470 44.510 80.050 44.680 ;
        RECT 75.530 44.030 75.950 44.240 ;
        RECT 76.420 44.030 76.840 44.240 ;
        RECT 77.650 44.070 79.110 44.240 ;
        RECT 75.600 43.970 75.860 44.030 ;
        RECT 76.510 43.970 76.770 44.030 ;
        RECT 74.020 43.190 74.190 43.900 ;
        RECT 71.990 42.750 72.250 42.840 ;
        RECT 72.900 42.750 73.160 42.840 ;
        RECT 69.670 42.540 71.090 42.710 ;
        RECT 71.900 42.540 72.320 42.750 ;
        RECT 72.830 42.540 73.250 42.750 ;
        RECT 68.730 42.100 70.310 42.270 ;
        RECT 71.520 42.150 71.690 42.480 ;
        RECT 65.560 41.330 65.730 41.660 ;
        RECT 66.970 41.540 68.550 41.710 ;
        RECT 64.030 41.060 64.450 41.270 ;
        RECT 64.920 41.060 65.340 41.270 ;
        RECT 66.150 41.100 67.610 41.270 ;
        RECT 64.100 41.000 64.360 41.060 ;
        RECT 65.010 41.000 65.270 41.060 ;
        RECT 66.610 41.040 66.900 41.100 ;
        RECT 68.130 40.930 68.550 41.270 ;
        RECT 68.810 41.230 68.980 42.100 ;
        RECT 69.360 41.230 69.530 41.920 ;
        RECT 73.500 41.880 73.670 42.570 ;
        RECT 74.040 41.710 74.210 42.580 ;
        RECT 74.480 42.540 74.900 42.820 ;
        RECT 76.120 42.710 76.290 43.280 ;
        RECT 77.770 43.190 77.940 44.070 ;
        RECT 78.110 44.010 78.400 44.070 ;
        RECT 79.630 43.900 80.050 44.240 ;
        RECT 80.310 44.200 80.480 45.070 ;
        RECT 80.860 44.200 81.030 44.890 ;
        RECT 85.000 44.850 85.170 45.540 ;
        RECT 85.540 44.680 85.710 45.550 ;
        RECT 85.980 45.510 86.400 45.790 ;
        RECT 87.620 45.680 87.790 46.010 ;
        RECT 89.240 45.720 89.500 45.810 ;
        RECT 90.150 45.720 90.410 45.810 ;
        RECT 86.920 45.510 88.340 45.680 ;
        RECT 89.150 45.510 89.570 45.720 ;
        RECT 90.080 45.510 90.500 45.720 ;
        RECT 85.980 45.070 87.560 45.240 ;
        RECT 88.770 45.120 88.940 45.450 ;
        RECT 82.810 44.300 82.980 44.630 ;
        RECT 84.220 44.510 85.800 44.680 ;
        RECT 81.280 44.030 81.700 44.240 ;
        RECT 82.170 44.030 82.590 44.240 ;
        RECT 83.400 44.070 84.860 44.240 ;
        RECT 81.350 43.970 81.610 44.030 ;
        RECT 82.260 43.970 82.520 44.030 ;
        RECT 79.770 43.190 79.940 43.900 ;
        RECT 77.740 42.750 78.000 42.840 ;
        RECT 78.650 42.750 78.910 42.840 ;
        RECT 75.420 42.540 76.840 42.710 ;
        RECT 77.650 42.540 78.070 42.750 ;
        RECT 78.580 42.540 79.000 42.750 ;
        RECT 74.480 42.100 76.060 42.270 ;
        RECT 77.270 42.150 77.440 42.480 ;
        RECT 71.310 41.330 71.480 41.660 ;
        RECT 72.720 41.540 74.300 41.710 ;
        RECT 69.780 41.060 70.200 41.270 ;
        RECT 70.670 41.060 71.090 41.270 ;
        RECT 71.900 41.100 73.360 41.270 ;
        RECT 69.850 41.000 70.110 41.060 ;
        RECT 70.760 41.000 71.020 41.060 ;
        RECT 72.360 41.040 72.650 41.100 ;
        RECT 73.880 40.930 74.300 41.270 ;
        RECT 74.560 41.230 74.730 42.100 ;
        RECT 75.110 41.230 75.280 41.920 ;
        RECT 79.250 41.880 79.420 42.570 ;
        RECT 79.790 41.710 79.960 42.580 ;
        RECT 80.230 42.540 80.650 42.820 ;
        RECT 81.870 42.710 82.040 43.280 ;
        RECT 83.520 43.190 83.690 44.070 ;
        RECT 83.860 44.010 84.150 44.070 ;
        RECT 85.380 43.900 85.800 44.240 ;
        RECT 86.060 44.200 86.230 45.070 ;
        RECT 86.610 44.200 86.780 44.890 ;
        RECT 90.750 44.850 90.920 45.540 ;
        RECT 91.290 44.680 91.460 45.550 ;
        RECT 91.730 45.510 92.150 45.790 ;
        RECT 93.370 45.680 93.540 46.010 ;
        RECT 92.670 45.510 94.090 45.680 ;
        RECT 91.730 45.070 93.310 45.240 ;
        RECT 88.560 44.300 88.730 44.630 ;
        RECT 89.970 44.510 91.550 44.680 ;
        RECT 87.030 44.030 87.450 44.240 ;
        RECT 87.920 44.030 88.340 44.240 ;
        RECT 89.150 44.070 90.610 44.240 ;
        RECT 87.100 43.970 87.360 44.030 ;
        RECT 88.010 43.970 88.270 44.030 ;
        RECT 85.520 43.190 85.690 43.900 ;
        RECT 83.490 42.750 83.750 42.840 ;
        RECT 84.400 42.750 84.660 42.840 ;
        RECT 81.170 42.540 82.590 42.710 ;
        RECT 83.400 42.540 83.820 42.750 ;
        RECT 84.330 42.540 84.750 42.750 ;
        RECT 80.230 42.100 81.810 42.270 ;
        RECT 83.020 42.150 83.190 42.480 ;
        RECT 77.060 41.330 77.230 41.660 ;
        RECT 78.470 41.540 80.050 41.710 ;
        RECT 75.530 41.060 75.950 41.270 ;
        RECT 76.420 41.060 76.840 41.270 ;
        RECT 77.650 41.100 79.110 41.270 ;
        RECT 75.600 41.000 75.860 41.060 ;
        RECT 76.510 41.000 76.770 41.060 ;
        RECT 78.110 41.040 78.400 41.100 ;
        RECT 79.630 40.930 80.050 41.270 ;
        RECT 80.310 41.230 80.480 42.100 ;
        RECT 80.860 41.230 81.030 41.920 ;
        RECT 85.000 41.880 85.170 42.570 ;
        RECT 85.540 41.710 85.710 42.580 ;
        RECT 85.980 42.540 86.400 42.820 ;
        RECT 87.620 42.710 87.790 43.280 ;
        RECT 89.270 43.190 89.440 44.070 ;
        RECT 89.610 44.010 89.900 44.070 ;
        RECT 91.130 43.900 91.550 44.240 ;
        RECT 91.810 44.200 91.980 45.070 ;
        RECT 92.360 44.200 92.530 44.890 ;
        RECT 94.310 44.300 94.480 44.630 ;
        RECT 92.780 44.030 93.200 44.240 ;
        RECT 93.670 44.030 94.090 44.240 ;
        RECT 92.850 43.970 93.110 44.030 ;
        RECT 93.760 43.970 94.020 44.030 ;
        RECT 91.270 43.190 91.440 43.900 ;
        RECT 94.230 43.280 94.400 43.550 ;
        RECT 93.370 43.110 94.400 43.280 ;
        RECT 89.240 42.750 89.500 42.840 ;
        RECT 90.150 42.750 90.410 42.840 ;
        RECT 86.920 42.540 88.340 42.710 ;
        RECT 89.150 42.540 89.570 42.750 ;
        RECT 90.080 42.540 90.500 42.750 ;
        RECT 85.980 42.100 87.560 42.270 ;
        RECT 88.770 42.150 88.940 42.480 ;
        RECT 82.810 41.330 82.980 41.660 ;
        RECT 84.220 41.540 85.800 41.710 ;
        RECT 81.280 41.060 81.700 41.270 ;
        RECT 82.170 41.060 82.590 41.270 ;
        RECT 83.400 41.100 84.860 41.270 ;
        RECT 81.350 41.000 81.610 41.060 ;
        RECT 82.260 41.000 82.520 41.060 ;
        RECT 83.860 41.040 84.150 41.100 ;
        RECT 85.380 40.930 85.800 41.270 ;
        RECT 86.060 41.230 86.230 42.100 ;
        RECT 86.610 41.230 86.780 41.920 ;
        RECT 90.750 41.880 90.920 42.570 ;
        RECT 91.290 41.710 91.460 42.580 ;
        RECT 91.730 42.540 92.150 42.820 ;
        RECT 93.370 42.710 93.540 43.110 ;
        RECT 92.670 42.540 94.090 42.710 ;
        RECT 91.730 42.100 93.310 42.270 ;
        RECT 88.560 41.330 88.730 41.660 ;
        RECT 89.970 41.540 91.550 41.710 ;
        RECT 87.030 41.060 87.450 41.270 ;
        RECT 87.920 41.060 88.340 41.270 ;
        RECT 89.150 41.100 90.610 41.270 ;
        RECT 87.100 41.000 87.360 41.060 ;
        RECT 88.010 41.000 88.270 41.060 ;
        RECT 89.610 41.040 89.900 41.100 ;
        RECT 91.130 40.930 91.550 41.270 ;
        RECT 91.810 41.230 91.980 42.100 ;
        RECT 92.360 41.230 92.530 41.920 ;
        RECT 94.310 41.330 94.480 41.660 ;
        RECT 92.780 41.060 93.200 41.270 ;
        RECT 93.670 41.060 94.090 41.270 ;
        RECT 92.850 41.000 93.110 41.060 ;
        RECT 93.760 41.000 94.020 41.060 ;
        RECT 2.990 40.340 3.250 40.430 ;
        RECT 3.900 40.340 4.160 40.430 ;
        RECT 2.900 40.130 3.320 40.340 ;
        RECT 3.830 40.130 4.250 40.340 ;
        RECT 2.520 39.740 2.690 40.070 ;
        RECT 4.500 39.470 4.670 40.160 ;
        RECT 5.040 39.300 5.210 40.170 ;
        RECT 5.480 40.130 5.900 40.410 ;
        RECT 7.120 40.300 7.290 40.630 ;
        RECT 8.740 40.340 9.000 40.430 ;
        RECT 9.650 40.340 9.910 40.430 ;
        RECT 6.420 40.130 7.840 40.300 ;
        RECT 8.650 40.130 9.070 40.340 ;
        RECT 9.580 40.130 10.000 40.340 ;
        RECT 5.480 39.690 7.060 39.860 ;
        RECT 8.270 39.740 8.440 40.070 ;
        RECT 3.720 39.130 5.300 39.300 ;
        RECT 2.900 38.690 4.360 38.860 ;
        RECT 3.360 38.630 3.650 38.690 ;
        RECT 4.880 38.520 5.300 38.860 ;
        RECT 5.560 38.820 5.730 39.690 ;
        RECT 6.110 38.820 6.280 39.510 ;
        RECT 10.250 39.470 10.420 40.160 ;
        RECT 10.790 39.300 10.960 40.170 ;
        RECT 11.230 40.130 11.650 40.410 ;
        RECT 12.870 40.300 13.040 40.630 ;
        RECT 14.490 40.340 14.750 40.430 ;
        RECT 15.400 40.340 15.660 40.430 ;
        RECT 12.170 40.130 13.590 40.300 ;
        RECT 14.400 40.130 14.820 40.340 ;
        RECT 15.330 40.130 15.750 40.340 ;
        RECT 11.230 39.690 12.810 39.860 ;
        RECT 14.020 39.740 14.190 40.070 ;
        RECT 8.060 38.920 8.230 39.250 ;
        RECT 9.470 39.130 11.050 39.300 ;
        RECT 6.530 38.650 6.950 38.860 ;
        RECT 7.420 38.650 7.840 38.860 ;
        RECT 8.650 38.690 10.110 38.860 ;
        RECT 6.600 38.590 6.860 38.650 ;
        RECT 7.510 38.590 7.770 38.650 ;
        RECT 9.110 38.630 9.400 38.690 ;
        RECT 10.630 38.520 11.050 38.860 ;
        RECT 11.310 38.820 11.480 39.690 ;
        RECT 11.860 38.820 12.030 39.510 ;
        RECT 16.000 39.470 16.170 40.160 ;
        RECT 16.540 39.300 16.710 40.170 ;
        RECT 16.980 40.130 17.400 40.410 ;
        RECT 18.620 40.300 18.790 40.630 ;
        RECT 20.240 40.340 20.500 40.430 ;
        RECT 21.150 40.340 21.410 40.430 ;
        RECT 17.920 40.130 19.340 40.300 ;
        RECT 20.150 40.130 20.570 40.340 ;
        RECT 21.080 40.130 21.500 40.340 ;
        RECT 16.980 39.690 18.560 39.860 ;
        RECT 19.770 39.740 19.940 40.070 ;
        RECT 13.810 38.920 13.980 39.250 ;
        RECT 15.220 39.130 16.800 39.300 ;
        RECT 12.280 38.650 12.700 38.860 ;
        RECT 13.170 38.650 13.590 38.860 ;
        RECT 14.400 38.690 15.860 38.860 ;
        RECT 12.350 38.590 12.610 38.650 ;
        RECT 13.260 38.590 13.520 38.650 ;
        RECT 14.860 38.630 15.150 38.690 ;
        RECT 16.380 38.520 16.800 38.860 ;
        RECT 17.060 38.820 17.230 39.690 ;
        RECT 17.610 38.820 17.780 39.510 ;
        RECT 21.750 39.470 21.920 40.160 ;
        RECT 22.290 39.300 22.460 40.170 ;
        RECT 22.730 40.130 23.150 40.410 ;
        RECT 24.370 40.300 24.540 40.630 ;
        RECT 25.990 40.340 26.250 40.430 ;
        RECT 26.900 40.340 27.160 40.430 ;
        RECT 23.670 40.130 25.090 40.300 ;
        RECT 25.900 40.130 26.320 40.340 ;
        RECT 26.830 40.130 27.250 40.340 ;
        RECT 22.730 39.690 24.310 39.860 ;
        RECT 25.520 39.740 25.690 40.070 ;
        RECT 19.560 38.920 19.730 39.250 ;
        RECT 20.970 39.130 22.550 39.300 ;
        RECT 18.030 38.650 18.450 38.860 ;
        RECT 18.920 38.650 19.340 38.860 ;
        RECT 20.150 38.690 21.610 38.860 ;
        RECT 18.100 38.590 18.360 38.650 ;
        RECT 19.010 38.590 19.270 38.650 ;
        RECT 20.610 38.630 20.900 38.690 ;
        RECT 22.130 38.520 22.550 38.860 ;
        RECT 22.810 38.820 22.980 39.690 ;
        RECT 23.360 38.820 23.530 39.510 ;
        RECT 27.500 39.470 27.670 40.160 ;
        RECT 28.040 39.300 28.210 40.170 ;
        RECT 28.480 40.130 28.900 40.410 ;
        RECT 30.120 40.300 30.290 40.630 ;
        RECT 31.740 40.340 32.000 40.430 ;
        RECT 32.650 40.340 32.910 40.430 ;
        RECT 29.420 40.130 30.840 40.300 ;
        RECT 31.650 40.130 32.070 40.340 ;
        RECT 32.580 40.130 33.000 40.340 ;
        RECT 28.480 39.690 30.060 39.860 ;
        RECT 31.270 39.740 31.440 40.070 ;
        RECT 25.310 38.920 25.480 39.250 ;
        RECT 26.720 39.130 28.300 39.300 ;
        RECT 23.780 38.650 24.200 38.860 ;
        RECT 24.670 38.650 25.090 38.860 ;
        RECT 25.900 38.690 27.360 38.860 ;
        RECT 23.850 38.590 24.110 38.650 ;
        RECT 24.760 38.590 25.020 38.650 ;
        RECT 26.360 38.630 26.650 38.690 ;
        RECT 27.880 38.520 28.300 38.860 ;
        RECT 28.560 38.820 28.730 39.690 ;
        RECT 29.110 38.820 29.280 39.510 ;
        RECT 33.250 39.470 33.420 40.160 ;
        RECT 33.790 39.300 33.960 40.170 ;
        RECT 34.230 40.130 34.650 40.410 ;
        RECT 35.870 40.300 36.040 40.630 ;
        RECT 37.490 40.340 37.750 40.430 ;
        RECT 38.400 40.340 38.660 40.430 ;
        RECT 35.170 40.130 36.590 40.300 ;
        RECT 37.400 40.130 37.820 40.340 ;
        RECT 38.330 40.130 38.750 40.340 ;
        RECT 34.230 39.690 35.810 39.860 ;
        RECT 37.020 39.740 37.190 40.070 ;
        RECT 31.060 38.920 31.230 39.250 ;
        RECT 32.470 39.130 34.050 39.300 ;
        RECT 29.530 38.650 29.950 38.860 ;
        RECT 30.420 38.650 30.840 38.860 ;
        RECT 31.650 38.690 33.110 38.860 ;
        RECT 29.600 38.590 29.860 38.650 ;
        RECT 30.510 38.590 30.770 38.650 ;
        RECT 32.110 38.630 32.400 38.690 ;
        RECT 33.630 38.520 34.050 38.860 ;
        RECT 34.310 38.820 34.480 39.690 ;
        RECT 34.860 38.820 35.030 39.510 ;
        RECT 39.000 39.470 39.170 40.160 ;
        RECT 39.540 39.300 39.710 40.170 ;
        RECT 39.980 40.130 40.400 40.410 ;
        RECT 41.620 40.300 41.790 40.630 ;
        RECT 43.240 40.340 43.500 40.430 ;
        RECT 44.150 40.340 44.410 40.430 ;
        RECT 40.920 40.130 42.340 40.300 ;
        RECT 43.150 40.130 43.570 40.340 ;
        RECT 44.080 40.130 44.500 40.340 ;
        RECT 39.980 39.690 41.560 39.860 ;
        RECT 42.770 39.740 42.940 40.070 ;
        RECT 36.810 38.920 36.980 39.250 ;
        RECT 38.220 39.130 39.800 39.300 ;
        RECT 35.280 38.650 35.700 38.860 ;
        RECT 36.170 38.650 36.590 38.860 ;
        RECT 37.400 38.690 38.860 38.860 ;
        RECT 35.350 38.590 35.610 38.650 ;
        RECT 36.260 38.590 36.520 38.650 ;
        RECT 37.860 38.630 38.150 38.690 ;
        RECT 39.380 38.520 39.800 38.860 ;
        RECT 40.060 38.820 40.230 39.690 ;
        RECT 40.610 38.820 40.780 39.510 ;
        RECT 44.750 39.470 44.920 40.160 ;
        RECT 45.290 39.300 45.460 40.170 ;
        RECT 45.730 40.130 46.150 40.410 ;
        RECT 47.370 40.300 47.540 40.630 ;
        RECT 48.990 40.340 49.250 40.430 ;
        RECT 49.900 40.340 50.160 40.430 ;
        RECT 46.670 40.130 48.090 40.300 ;
        RECT 48.900 40.130 49.320 40.340 ;
        RECT 49.830 40.130 50.250 40.340 ;
        RECT 45.730 39.690 47.310 39.860 ;
        RECT 48.520 39.740 48.690 40.070 ;
        RECT 42.560 38.920 42.730 39.250 ;
        RECT 43.970 39.130 45.550 39.300 ;
        RECT 41.030 38.650 41.450 38.860 ;
        RECT 41.920 38.650 42.340 38.860 ;
        RECT 43.150 38.690 44.610 38.860 ;
        RECT 41.100 38.590 41.360 38.650 ;
        RECT 42.010 38.590 42.270 38.650 ;
        RECT 43.610 38.630 43.900 38.690 ;
        RECT 45.130 38.520 45.550 38.860 ;
        RECT 45.810 38.820 45.980 39.690 ;
        RECT 46.360 38.820 46.530 39.510 ;
        RECT 50.500 39.470 50.670 40.160 ;
        RECT 51.040 39.300 51.210 40.170 ;
        RECT 51.480 40.130 51.900 40.410 ;
        RECT 53.120 40.300 53.290 40.630 ;
        RECT 54.740 40.340 55.000 40.430 ;
        RECT 55.650 40.340 55.910 40.430 ;
        RECT 52.420 40.130 53.840 40.300 ;
        RECT 54.650 40.130 55.070 40.340 ;
        RECT 55.580 40.130 56.000 40.340 ;
        RECT 51.480 39.690 53.060 39.860 ;
        RECT 54.270 39.740 54.440 40.070 ;
        RECT 48.310 38.920 48.480 39.250 ;
        RECT 49.720 39.130 51.300 39.300 ;
        RECT 46.780 38.650 47.200 38.860 ;
        RECT 47.670 38.650 48.090 38.860 ;
        RECT 48.900 38.690 50.360 38.860 ;
        RECT 46.850 38.590 47.110 38.650 ;
        RECT 47.760 38.590 48.020 38.650 ;
        RECT 49.360 38.630 49.650 38.690 ;
        RECT 50.880 38.520 51.300 38.860 ;
        RECT 51.560 38.820 51.730 39.690 ;
        RECT 52.110 38.820 52.280 39.510 ;
        RECT 56.250 39.470 56.420 40.160 ;
        RECT 56.790 39.300 56.960 40.170 ;
        RECT 57.230 40.130 57.650 40.410 ;
        RECT 58.870 40.300 59.040 40.630 ;
        RECT 60.490 40.340 60.750 40.430 ;
        RECT 61.400 40.340 61.660 40.430 ;
        RECT 58.170 40.130 59.590 40.300 ;
        RECT 60.400 40.130 60.820 40.340 ;
        RECT 61.330 40.130 61.750 40.340 ;
        RECT 57.230 39.690 58.810 39.860 ;
        RECT 60.020 39.740 60.190 40.070 ;
        RECT 54.060 38.920 54.230 39.250 ;
        RECT 55.470 39.130 57.050 39.300 ;
        RECT 52.530 38.650 52.950 38.860 ;
        RECT 53.420 38.650 53.840 38.860 ;
        RECT 54.650 38.690 56.110 38.860 ;
        RECT 52.600 38.590 52.860 38.650 ;
        RECT 53.510 38.590 53.770 38.650 ;
        RECT 55.110 38.630 55.400 38.690 ;
        RECT 56.630 38.520 57.050 38.860 ;
        RECT 57.310 38.820 57.480 39.690 ;
        RECT 57.860 38.820 58.030 39.510 ;
        RECT 62.000 39.470 62.170 40.160 ;
        RECT 62.540 39.300 62.710 40.170 ;
        RECT 62.980 40.130 63.400 40.410 ;
        RECT 64.620 40.300 64.790 40.630 ;
        RECT 66.240 40.340 66.500 40.430 ;
        RECT 67.150 40.340 67.410 40.430 ;
        RECT 63.920 40.130 65.340 40.300 ;
        RECT 66.150 40.130 66.570 40.340 ;
        RECT 67.080 40.130 67.500 40.340 ;
        RECT 62.980 39.690 64.560 39.860 ;
        RECT 65.770 39.740 65.940 40.070 ;
        RECT 59.810 38.920 59.980 39.250 ;
        RECT 61.220 39.130 62.800 39.300 ;
        RECT 58.280 38.650 58.700 38.860 ;
        RECT 59.170 38.650 59.590 38.860 ;
        RECT 60.400 38.690 61.860 38.860 ;
        RECT 58.350 38.590 58.610 38.650 ;
        RECT 59.260 38.590 59.520 38.650 ;
        RECT 60.860 38.630 61.150 38.690 ;
        RECT 62.380 38.520 62.800 38.860 ;
        RECT 63.060 38.820 63.230 39.690 ;
        RECT 63.610 38.820 63.780 39.510 ;
        RECT 67.750 39.470 67.920 40.160 ;
        RECT 68.290 39.300 68.460 40.170 ;
        RECT 68.730 40.130 69.150 40.410 ;
        RECT 70.370 40.300 70.540 40.630 ;
        RECT 71.990 40.340 72.250 40.430 ;
        RECT 72.900 40.340 73.160 40.430 ;
        RECT 69.670 40.130 71.090 40.300 ;
        RECT 71.900 40.130 72.320 40.340 ;
        RECT 72.830 40.130 73.250 40.340 ;
        RECT 68.730 39.690 70.310 39.860 ;
        RECT 71.520 39.740 71.690 40.070 ;
        RECT 65.560 38.920 65.730 39.250 ;
        RECT 66.970 39.130 68.550 39.300 ;
        RECT 64.030 38.650 64.450 38.860 ;
        RECT 64.920 38.650 65.340 38.860 ;
        RECT 66.150 38.690 67.610 38.860 ;
        RECT 64.100 38.590 64.360 38.650 ;
        RECT 65.010 38.590 65.270 38.650 ;
        RECT 66.610 38.630 66.900 38.690 ;
        RECT 68.130 38.520 68.550 38.860 ;
        RECT 68.810 38.820 68.980 39.690 ;
        RECT 69.360 38.820 69.530 39.510 ;
        RECT 73.500 39.470 73.670 40.160 ;
        RECT 74.040 39.300 74.210 40.170 ;
        RECT 74.480 40.130 74.900 40.410 ;
        RECT 76.120 40.300 76.290 40.630 ;
        RECT 77.740 40.340 78.000 40.430 ;
        RECT 78.650 40.340 78.910 40.430 ;
        RECT 75.420 40.130 76.840 40.300 ;
        RECT 77.650 40.130 78.070 40.340 ;
        RECT 78.580 40.130 79.000 40.340 ;
        RECT 74.480 39.690 76.060 39.860 ;
        RECT 77.270 39.740 77.440 40.070 ;
        RECT 71.310 38.920 71.480 39.250 ;
        RECT 72.720 39.130 74.300 39.300 ;
        RECT 69.780 38.650 70.200 38.860 ;
        RECT 70.670 38.650 71.090 38.860 ;
        RECT 71.900 38.690 73.360 38.860 ;
        RECT 69.850 38.590 70.110 38.650 ;
        RECT 70.760 38.590 71.020 38.650 ;
        RECT 72.360 38.630 72.650 38.690 ;
        RECT 73.880 38.520 74.300 38.860 ;
        RECT 74.560 38.820 74.730 39.690 ;
        RECT 75.110 38.820 75.280 39.510 ;
        RECT 79.250 39.470 79.420 40.160 ;
        RECT 79.790 39.300 79.960 40.170 ;
        RECT 80.230 40.130 80.650 40.410 ;
        RECT 81.870 40.300 82.040 40.630 ;
        RECT 83.490 40.340 83.750 40.430 ;
        RECT 84.400 40.340 84.660 40.430 ;
        RECT 81.170 40.130 82.590 40.300 ;
        RECT 83.400 40.130 83.820 40.340 ;
        RECT 84.330 40.130 84.750 40.340 ;
        RECT 80.230 39.690 81.810 39.860 ;
        RECT 83.020 39.740 83.190 40.070 ;
        RECT 77.060 38.920 77.230 39.250 ;
        RECT 78.470 39.130 80.050 39.300 ;
        RECT 75.530 38.650 75.950 38.860 ;
        RECT 76.420 38.650 76.840 38.860 ;
        RECT 77.650 38.690 79.110 38.860 ;
        RECT 75.600 38.590 75.860 38.650 ;
        RECT 76.510 38.590 76.770 38.650 ;
        RECT 78.110 38.630 78.400 38.690 ;
        RECT 79.630 38.520 80.050 38.860 ;
        RECT 80.310 38.820 80.480 39.690 ;
        RECT 80.860 38.820 81.030 39.510 ;
        RECT 85.000 39.470 85.170 40.160 ;
        RECT 85.540 39.300 85.710 40.170 ;
        RECT 85.980 40.130 86.400 40.410 ;
        RECT 87.620 40.300 87.790 40.630 ;
        RECT 89.240 40.340 89.500 40.430 ;
        RECT 90.150 40.340 90.410 40.430 ;
        RECT 86.920 40.130 88.340 40.300 ;
        RECT 89.150 40.130 89.570 40.340 ;
        RECT 90.080 40.130 90.500 40.340 ;
        RECT 85.980 39.690 87.560 39.860 ;
        RECT 88.770 39.740 88.940 40.070 ;
        RECT 82.810 38.920 82.980 39.250 ;
        RECT 84.220 39.130 85.800 39.300 ;
        RECT 81.280 38.650 81.700 38.860 ;
        RECT 82.170 38.650 82.590 38.860 ;
        RECT 83.400 38.690 84.860 38.860 ;
        RECT 81.350 38.590 81.610 38.650 ;
        RECT 82.260 38.590 82.520 38.650 ;
        RECT 83.860 38.630 84.150 38.690 ;
        RECT 85.380 38.520 85.800 38.860 ;
        RECT 86.060 38.820 86.230 39.690 ;
        RECT 86.610 38.820 86.780 39.510 ;
        RECT 90.750 39.470 90.920 40.160 ;
        RECT 91.290 39.300 91.460 40.170 ;
        RECT 91.730 40.130 92.150 40.410 ;
        RECT 93.370 40.300 93.540 40.630 ;
        RECT 92.670 40.130 94.090 40.300 ;
        RECT 91.730 39.690 93.310 39.860 ;
        RECT 88.560 38.920 88.730 39.250 ;
        RECT 89.970 39.130 91.550 39.300 ;
        RECT 87.030 38.650 87.450 38.860 ;
        RECT 87.920 38.650 88.340 38.860 ;
        RECT 89.150 38.690 90.610 38.860 ;
        RECT 87.100 38.590 87.360 38.650 ;
        RECT 88.010 38.590 88.270 38.650 ;
        RECT 89.610 38.630 89.900 38.690 ;
        RECT 91.130 38.520 91.550 38.860 ;
        RECT 91.810 38.820 91.980 39.690 ;
        RECT 92.360 38.820 92.530 39.510 ;
        RECT 94.310 38.920 94.480 39.250 ;
        RECT 92.780 38.650 93.200 38.860 ;
        RECT 93.670 38.650 94.090 38.860 ;
        RECT 92.850 38.590 93.110 38.650 ;
        RECT 93.760 38.590 94.020 38.650 ;
        RECT 2.990 37.930 3.250 38.020 ;
        RECT 3.900 37.930 4.160 38.020 ;
        RECT 2.900 37.720 3.320 37.930 ;
        RECT 3.830 37.720 4.250 37.930 ;
        RECT 2.520 37.330 2.690 37.660 ;
        RECT 4.500 37.060 4.670 37.750 ;
        RECT 5.040 36.890 5.210 37.760 ;
        RECT 5.480 37.720 5.900 38.000 ;
        RECT 7.120 37.890 7.290 38.220 ;
        RECT 8.740 37.930 9.000 38.020 ;
        RECT 9.650 37.930 9.910 38.020 ;
        RECT 6.420 37.720 7.840 37.890 ;
        RECT 8.650 37.720 9.070 37.930 ;
        RECT 9.580 37.720 10.000 37.930 ;
        RECT 5.480 37.280 7.060 37.450 ;
        RECT 8.270 37.330 8.440 37.660 ;
        RECT 3.720 36.720 5.300 36.890 ;
        RECT 2.900 36.280 4.360 36.450 ;
        RECT 3.360 36.220 3.650 36.280 ;
        RECT 4.880 36.110 5.300 36.450 ;
        RECT 5.560 36.410 5.730 37.280 ;
        RECT 6.110 36.410 6.280 37.100 ;
        RECT 10.250 37.060 10.420 37.750 ;
        RECT 10.790 36.890 10.960 37.760 ;
        RECT 11.230 37.720 11.650 38.000 ;
        RECT 12.870 37.890 13.040 38.220 ;
        RECT 14.490 37.930 14.750 38.020 ;
        RECT 15.400 37.930 15.660 38.020 ;
        RECT 12.170 37.720 13.590 37.890 ;
        RECT 14.400 37.720 14.820 37.930 ;
        RECT 15.330 37.720 15.750 37.930 ;
        RECT 11.230 37.280 12.810 37.450 ;
        RECT 14.020 37.330 14.190 37.660 ;
        RECT 8.060 36.510 8.230 36.840 ;
        RECT 9.470 36.720 11.050 36.890 ;
        RECT 6.530 36.240 6.950 36.450 ;
        RECT 7.420 36.240 7.840 36.450 ;
        RECT 8.650 36.280 10.110 36.450 ;
        RECT 6.600 36.180 6.860 36.240 ;
        RECT 7.510 36.180 7.770 36.240 ;
        RECT 9.110 36.220 9.400 36.280 ;
        RECT 10.630 36.110 11.050 36.450 ;
        RECT 11.310 36.410 11.480 37.280 ;
        RECT 11.860 36.410 12.030 37.100 ;
        RECT 16.000 37.060 16.170 37.750 ;
        RECT 16.540 36.890 16.710 37.760 ;
        RECT 16.980 37.720 17.400 38.000 ;
        RECT 18.620 37.890 18.790 38.220 ;
        RECT 20.240 37.930 20.500 38.020 ;
        RECT 21.150 37.930 21.410 38.020 ;
        RECT 17.920 37.720 19.340 37.890 ;
        RECT 20.150 37.720 20.570 37.930 ;
        RECT 21.080 37.720 21.500 37.930 ;
        RECT 16.980 37.280 18.560 37.450 ;
        RECT 19.770 37.330 19.940 37.660 ;
        RECT 13.810 36.510 13.980 36.840 ;
        RECT 15.220 36.720 16.800 36.890 ;
        RECT 12.280 36.240 12.700 36.450 ;
        RECT 13.170 36.240 13.590 36.450 ;
        RECT 14.400 36.280 15.860 36.450 ;
        RECT 12.350 36.180 12.610 36.240 ;
        RECT 13.260 36.180 13.520 36.240 ;
        RECT 14.860 36.220 15.150 36.280 ;
        RECT 16.380 36.110 16.800 36.450 ;
        RECT 17.060 36.410 17.230 37.280 ;
        RECT 17.610 36.410 17.780 37.100 ;
        RECT 21.750 37.060 21.920 37.750 ;
        RECT 22.290 36.890 22.460 37.760 ;
        RECT 22.730 37.720 23.150 38.000 ;
        RECT 24.370 37.890 24.540 38.220 ;
        RECT 25.990 37.930 26.250 38.020 ;
        RECT 26.900 37.930 27.160 38.020 ;
        RECT 23.670 37.720 25.090 37.890 ;
        RECT 25.900 37.720 26.320 37.930 ;
        RECT 26.830 37.720 27.250 37.930 ;
        RECT 22.730 37.280 24.310 37.450 ;
        RECT 25.520 37.330 25.690 37.660 ;
        RECT 19.560 36.510 19.730 36.840 ;
        RECT 20.970 36.720 22.550 36.890 ;
        RECT 18.030 36.240 18.450 36.450 ;
        RECT 18.920 36.240 19.340 36.450 ;
        RECT 20.150 36.280 21.610 36.450 ;
        RECT 18.100 36.180 18.360 36.240 ;
        RECT 19.010 36.180 19.270 36.240 ;
        RECT 20.610 36.220 20.900 36.280 ;
        RECT 22.130 36.110 22.550 36.450 ;
        RECT 22.810 36.410 22.980 37.280 ;
        RECT 23.360 36.410 23.530 37.100 ;
        RECT 27.500 37.060 27.670 37.750 ;
        RECT 28.040 36.890 28.210 37.760 ;
        RECT 28.480 37.720 28.900 38.000 ;
        RECT 30.120 37.890 30.290 38.220 ;
        RECT 31.740 37.930 32.000 38.020 ;
        RECT 32.650 37.930 32.910 38.020 ;
        RECT 29.420 37.720 30.840 37.890 ;
        RECT 31.650 37.720 32.070 37.930 ;
        RECT 32.580 37.720 33.000 37.930 ;
        RECT 28.480 37.280 30.060 37.450 ;
        RECT 31.270 37.330 31.440 37.660 ;
        RECT 25.310 36.510 25.480 36.840 ;
        RECT 26.720 36.720 28.300 36.890 ;
        RECT 23.780 36.240 24.200 36.450 ;
        RECT 24.670 36.240 25.090 36.450 ;
        RECT 25.900 36.280 27.360 36.450 ;
        RECT 23.850 36.180 24.110 36.240 ;
        RECT 24.760 36.180 25.020 36.240 ;
        RECT 26.360 36.220 26.650 36.280 ;
        RECT 27.880 36.110 28.300 36.450 ;
        RECT 28.560 36.410 28.730 37.280 ;
        RECT 29.110 36.410 29.280 37.100 ;
        RECT 33.250 37.060 33.420 37.750 ;
        RECT 33.790 36.890 33.960 37.760 ;
        RECT 34.230 37.720 34.650 38.000 ;
        RECT 35.870 37.890 36.040 38.220 ;
        RECT 37.490 37.930 37.750 38.020 ;
        RECT 38.400 37.930 38.660 38.020 ;
        RECT 35.170 37.720 36.590 37.890 ;
        RECT 37.400 37.720 37.820 37.930 ;
        RECT 38.330 37.720 38.750 37.930 ;
        RECT 34.230 37.280 35.810 37.450 ;
        RECT 37.020 37.330 37.190 37.660 ;
        RECT 31.060 36.510 31.230 36.840 ;
        RECT 32.470 36.720 34.050 36.890 ;
        RECT 29.530 36.240 29.950 36.450 ;
        RECT 30.420 36.240 30.840 36.450 ;
        RECT 31.650 36.280 33.110 36.450 ;
        RECT 29.600 36.180 29.860 36.240 ;
        RECT 30.510 36.180 30.770 36.240 ;
        RECT 32.110 36.220 32.400 36.280 ;
        RECT 33.630 36.110 34.050 36.450 ;
        RECT 34.310 36.410 34.480 37.280 ;
        RECT 34.860 36.410 35.030 37.100 ;
        RECT 39.000 37.060 39.170 37.750 ;
        RECT 39.540 36.890 39.710 37.760 ;
        RECT 39.980 37.720 40.400 38.000 ;
        RECT 41.620 37.890 41.790 38.220 ;
        RECT 43.240 37.930 43.500 38.020 ;
        RECT 44.150 37.930 44.410 38.020 ;
        RECT 40.920 37.720 42.340 37.890 ;
        RECT 43.150 37.720 43.570 37.930 ;
        RECT 44.080 37.720 44.500 37.930 ;
        RECT 39.980 37.280 41.560 37.450 ;
        RECT 42.770 37.330 42.940 37.660 ;
        RECT 36.810 36.510 36.980 36.840 ;
        RECT 38.220 36.720 39.800 36.890 ;
        RECT 35.280 36.240 35.700 36.450 ;
        RECT 36.170 36.240 36.590 36.450 ;
        RECT 37.400 36.280 38.860 36.450 ;
        RECT 35.350 36.180 35.610 36.240 ;
        RECT 36.260 36.180 36.520 36.240 ;
        RECT 37.860 36.220 38.150 36.280 ;
        RECT 39.380 36.110 39.800 36.450 ;
        RECT 40.060 36.410 40.230 37.280 ;
        RECT 40.610 36.410 40.780 37.100 ;
        RECT 44.750 37.060 44.920 37.750 ;
        RECT 45.290 36.890 45.460 37.760 ;
        RECT 45.730 37.720 46.150 38.000 ;
        RECT 47.370 37.890 47.540 38.220 ;
        RECT 48.990 37.930 49.250 38.020 ;
        RECT 49.900 37.930 50.160 38.020 ;
        RECT 46.670 37.720 48.090 37.890 ;
        RECT 48.900 37.720 49.320 37.930 ;
        RECT 49.830 37.720 50.250 37.930 ;
        RECT 45.730 37.280 47.310 37.450 ;
        RECT 48.520 37.330 48.690 37.660 ;
        RECT 42.560 36.510 42.730 36.840 ;
        RECT 43.970 36.720 45.550 36.890 ;
        RECT 41.030 36.240 41.450 36.450 ;
        RECT 41.920 36.240 42.340 36.450 ;
        RECT 43.150 36.280 44.610 36.450 ;
        RECT 41.100 36.180 41.360 36.240 ;
        RECT 42.010 36.180 42.270 36.240 ;
        RECT 43.610 36.220 43.900 36.280 ;
        RECT 45.130 36.110 45.550 36.450 ;
        RECT 45.810 36.410 45.980 37.280 ;
        RECT 46.360 36.410 46.530 37.100 ;
        RECT 50.500 37.060 50.670 37.750 ;
        RECT 51.040 36.890 51.210 37.760 ;
        RECT 51.480 37.720 51.900 38.000 ;
        RECT 53.120 37.890 53.290 38.220 ;
        RECT 54.740 37.930 55.000 38.020 ;
        RECT 55.650 37.930 55.910 38.020 ;
        RECT 52.420 37.720 53.840 37.890 ;
        RECT 54.650 37.720 55.070 37.930 ;
        RECT 55.580 37.720 56.000 37.930 ;
        RECT 51.480 37.280 53.060 37.450 ;
        RECT 54.270 37.330 54.440 37.660 ;
        RECT 48.310 36.510 48.480 36.840 ;
        RECT 49.720 36.720 51.300 36.890 ;
        RECT 46.780 36.240 47.200 36.450 ;
        RECT 47.670 36.240 48.090 36.450 ;
        RECT 48.900 36.280 50.360 36.450 ;
        RECT 46.850 36.180 47.110 36.240 ;
        RECT 47.760 36.180 48.020 36.240 ;
        RECT 49.360 36.220 49.650 36.280 ;
        RECT 50.880 36.110 51.300 36.450 ;
        RECT 51.560 36.410 51.730 37.280 ;
        RECT 52.110 36.410 52.280 37.100 ;
        RECT 56.250 37.060 56.420 37.750 ;
        RECT 56.790 36.890 56.960 37.760 ;
        RECT 57.230 37.720 57.650 38.000 ;
        RECT 58.870 37.890 59.040 38.220 ;
        RECT 60.490 37.930 60.750 38.020 ;
        RECT 61.400 37.930 61.660 38.020 ;
        RECT 58.170 37.720 59.590 37.890 ;
        RECT 60.400 37.720 60.820 37.930 ;
        RECT 61.330 37.720 61.750 37.930 ;
        RECT 57.230 37.280 58.810 37.450 ;
        RECT 60.020 37.330 60.190 37.660 ;
        RECT 54.060 36.510 54.230 36.840 ;
        RECT 55.470 36.720 57.050 36.890 ;
        RECT 52.530 36.240 52.950 36.450 ;
        RECT 53.420 36.240 53.840 36.450 ;
        RECT 54.650 36.280 56.110 36.450 ;
        RECT 52.600 36.180 52.860 36.240 ;
        RECT 53.510 36.180 53.770 36.240 ;
        RECT 55.110 36.220 55.400 36.280 ;
        RECT 56.630 36.110 57.050 36.450 ;
        RECT 57.310 36.410 57.480 37.280 ;
        RECT 57.860 36.410 58.030 37.100 ;
        RECT 62.000 37.060 62.170 37.750 ;
        RECT 62.540 36.890 62.710 37.760 ;
        RECT 62.980 37.720 63.400 38.000 ;
        RECT 64.620 37.890 64.790 38.220 ;
        RECT 66.240 37.930 66.500 38.020 ;
        RECT 67.150 37.930 67.410 38.020 ;
        RECT 63.920 37.720 65.340 37.890 ;
        RECT 66.150 37.720 66.570 37.930 ;
        RECT 67.080 37.720 67.500 37.930 ;
        RECT 62.980 37.280 64.560 37.450 ;
        RECT 65.770 37.330 65.940 37.660 ;
        RECT 59.810 36.510 59.980 36.840 ;
        RECT 61.220 36.720 62.800 36.890 ;
        RECT 58.280 36.240 58.700 36.450 ;
        RECT 59.170 36.240 59.590 36.450 ;
        RECT 60.400 36.280 61.860 36.450 ;
        RECT 58.350 36.180 58.610 36.240 ;
        RECT 59.260 36.180 59.520 36.240 ;
        RECT 60.860 36.220 61.150 36.280 ;
        RECT 62.380 36.110 62.800 36.450 ;
        RECT 63.060 36.410 63.230 37.280 ;
        RECT 63.610 36.410 63.780 37.100 ;
        RECT 67.750 37.060 67.920 37.750 ;
        RECT 68.290 36.890 68.460 37.760 ;
        RECT 68.730 37.720 69.150 38.000 ;
        RECT 70.370 37.890 70.540 38.220 ;
        RECT 71.990 37.930 72.250 38.020 ;
        RECT 72.900 37.930 73.160 38.020 ;
        RECT 69.670 37.720 71.090 37.890 ;
        RECT 71.900 37.720 72.320 37.930 ;
        RECT 72.830 37.720 73.250 37.930 ;
        RECT 68.730 37.280 70.310 37.450 ;
        RECT 71.520 37.330 71.690 37.660 ;
        RECT 65.560 36.510 65.730 36.840 ;
        RECT 66.970 36.720 68.550 36.890 ;
        RECT 64.030 36.240 64.450 36.450 ;
        RECT 64.920 36.240 65.340 36.450 ;
        RECT 66.150 36.280 67.610 36.450 ;
        RECT 64.100 36.180 64.360 36.240 ;
        RECT 65.010 36.180 65.270 36.240 ;
        RECT 66.610 36.220 66.900 36.280 ;
        RECT 68.130 36.110 68.550 36.450 ;
        RECT 68.810 36.410 68.980 37.280 ;
        RECT 69.360 36.410 69.530 37.100 ;
        RECT 73.500 37.060 73.670 37.750 ;
        RECT 74.040 36.890 74.210 37.760 ;
        RECT 74.480 37.720 74.900 38.000 ;
        RECT 76.120 37.890 76.290 38.220 ;
        RECT 77.740 37.930 78.000 38.020 ;
        RECT 78.650 37.930 78.910 38.020 ;
        RECT 75.420 37.720 76.840 37.890 ;
        RECT 77.650 37.720 78.070 37.930 ;
        RECT 78.580 37.720 79.000 37.930 ;
        RECT 74.480 37.280 76.060 37.450 ;
        RECT 77.270 37.330 77.440 37.660 ;
        RECT 71.310 36.510 71.480 36.840 ;
        RECT 72.720 36.720 74.300 36.890 ;
        RECT 69.780 36.240 70.200 36.450 ;
        RECT 70.670 36.240 71.090 36.450 ;
        RECT 71.900 36.280 73.360 36.450 ;
        RECT 69.850 36.180 70.110 36.240 ;
        RECT 70.760 36.180 71.020 36.240 ;
        RECT 72.360 36.220 72.650 36.280 ;
        RECT 73.880 36.110 74.300 36.450 ;
        RECT 74.560 36.410 74.730 37.280 ;
        RECT 75.110 36.410 75.280 37.100 ;
        RECT 79.250 37.060 79.420 37.750 ;
        RECT 79.790 36.890 79.960 37.760 ;
        RECT 80.230 37.720 80.650 38.000 ;
        RECT 81.870 37.890 82.040 38.220 ;
        RECT 83.490 37.930 83.750 38.020 ;
        RECT 84.400 37.930 84.660 38.020 ;
        RECT 81.170 37.720 82.590 37.890 ;
        RECT 83.400 37.720 83.820 37.930 ;
        RECT 84.330 37.720 84.750 37.930 ;
        RECT 80.230 37.280 81.810 37.450 ;
        RECT 83.020 37.330 83.190 37.660 ;
        RECT 77.060 36.510 77.230 36.840 ;
        RECT 78.470 36.720 80.050 36.890 ;
        RECT 75.530 36.240 75.950 36.450 ;
        RECT 76.420 36.240 76.840 36.450 ;
        RECT 77.650 36.280 79.110 36.450 ;
        RECT 75.600 36.180 75.860 36.240 ;
        RECT 76.510 36.180 76.770 36.240 ;
        RECT 78.110 36.220 78.400 36.280 ;
        RECT 79.630 36.110 80.050 36.450 ;
        RECT 80.310 36.410 80.480 37.280 ;
        RECT 80.860 36.410 81.030 37.100 ;
        RECT 85.000 37.060 85.170 37.750 ;
        RECT 85.540 36.890 85.710 37.760 ;
        RECT 85.980 37.720 86.400 38.000 ;
        RECT 87.620 37.890 87.790 38.220 ;
        RECT 89.240 37.930 89.500 38.020 ;
        RECT 90.150 37.930 90.410 38.020 ;
        RECT 86.920 37.720 88.340 37.890 ;
        RECT 89.150 37.720 89.570 37.930 ;
        RECT 90.080 37.720 90.500 37.930 ;
        RECT 85.980 37.280 87.560 37.450 ;
        RECT 88.770 37.330 88.940 37.660 ;
        RECT 82.810 36.510 82.980 36.840 ;
        RECT 84.220 36.720 85.800 36.890 ;
        RECT 81.280 36.240 81.700 36.450 ;
        RECT 82.170 36.240 82.590 36.450 ;
        RECT 83.400 36.280 84.860 36.450 ;
        RECT 81.350 36.180 81.610 36.240 ;
        RECT 82.260 36.180 82.520 36.240 ;
        RECT 83.860 36.220 84.150 36.280 ;
        RECT 85.380 36.110 85.800 36.450 ;
        RECT 86.060 36.410 86.230 37.280 ;
        RECT 86.610 36.410 86.780 37.100 ;
        RECT 90.750 37.060 90.920 37.750 ;
        RECT 91.290 36.890 91.460 37.760 ;
        RECT 91.730 37.720 92.150 38.000 ;
        RECT 93.370 37.890 93.540 38.220 ;
        RECT 92.670 37.720 94.090 37.890 ;
        RECT 91.730 37.280 93.310 37.450 ;
        RECT 88.560 36.510 88.730 36.840 ;
        RECT 89.970 36.720 91.550 36.890 ;
        RECT 87.030 36.240 87.450 36.450 ;
        RECT 87.920 36.240 88.340 36.450 ;
        RECT 89.150 36.280 90.610 36.450 ;
        RECT 87.100 36.180 87.360 36.240 ;
        RECT 88.010 36.180 88.270 36.240 ;
        RECT 89.610 36.220 89.900 36.280 ;
        RECT 91.130 36.110 91.550 36.450 ;
        RECT 91.810 36.410 91.980 37.280 ;
        RECT 92.360 36.410 92.530 37.100 ;
        RECT 94.310 36.510 94.480 36.840 ;
        RECT 92.780 36.240 93.200 36.450 ;
        RECT 93.670 36.240 94.090 36.450 ;
        RECT 92.850 36.180 93.110 36.240 ;
        RECT 93.760 36.180 94.020 36.240 ;
        RECT 2.990 35.520 3.250 35.610 ;
        RECT 3.900 35.520 4.160 35.610 ;
        RECT 2.900 35.310 3.320 35.520 ;
        RECT 3.830 35.310 4.250 35.520 ;
        RECT 2.520 34.920 2.690 35.250 ;
        RECT 4.500 34.650 4.670 35.340 ;
        RECT 5.040 34.480 5.210 35.350 ;
        RECT 5.480 35.310 5.900 35.590 ;
        RECT 7.120 35.480 7.290 35.810 ;
        RECT 8.740 35.520 9.000 35.610 ;
        RECT 9.650 35.520 9.910 35.610 ;
        RECT 6.420 35.310 7.840 35.480 ;
        RECT 8.650 35.310 9.070 35.520 ;
        RECT 9.580 35.310 10.000 35.520 ;
        RECT 5.480 34.870 7.060 35.040 ;
        RECT 8.270 34.920 8.440 35.250 ;
        RECT 3.720 34.310 5.300 34.480 ;
        RECT 2.900 33.870 4.360 34.040 ;
        RECT 3.360 33.810 3.650 33.870 ;
        RECT 4.880 33.700 5.300 34.040 ;
        RECT 5.560 34.000 5.730 34.870 ;
        RECT 6.110 34.000 6.280 34.690 ;
        RECT 10.250 34.650 10.420 35.340 ;
        RECT 10.790 34.480 10.960 35.350 ;
        RECT 11.230 35.310 11.650 35.590 ;
        RECT 12.870 35.480 13.040 35.810 ;
        RECT 14.490 35.520 14.750 35.610 ;
        RECT 15.400 35.520 15.660 35.610 ;
        RECT 12.170 35.310 13.590 35.480 ;
        RECT 14.400 35.310 14.820 35.520 ;
        RECT 15.330 35.310 15.750 35.520 ;
        RECT 11.230 34.870 12.810 35.040 ;
        RECT 14.020 34.920 14.190 35.250 ;
        RECT 8.060 34.100 8.230 34.430 ;
        RECT 9.470 34.310 11.050 34.480 ;
        RECT 6.530 33.830 6.950 34.040 ;
        RECT 7.420 33.830 7.840 34.040 ;
        RECT 8.650 33.870 10.110 34.040 ;
        RECT 6.600 33.770 6.860 33.830 ;
        RECT 7.510 33.770 7.770 33.830 ;
        RECT 9.110 33.810 9.400 33.870 ;
        RECT 10.630 33.700 11.050 34.040 ;
        RECT 11.310 34.000 11.480 34.870 ;
        RECT 11.860 34.000 12.030 34.690 ;
        RECT 16.000 34.650 16.170 35.340 ;
        RECT 16.540 34.480 16.710 35.350 ;
        RECT 16.980 35.310 17.400 35.590 ;
        RECT 18.620 35.480 18.790 35.810 ;
        RECT 20.240 35.520 20.500 35.610 ;
        RECT 21.150 35.520 21.410 35.610 ;
        RECT 17.920 35.310 19.340 35.480 ;
        RECT 20.150 35.310 20.570 35.520 ;
        RECT 21.080 35.310 21.500 35.520 ;
        RECT 16.980 34.870 18.560 35.040 ;
        RECT 19.770 34.920 19.940 35.250 ;
        RECT 13.810 34.100 13.980 34.430 ;
        RECT 15.220 34.310 16.800 34.480 ;
        RECT 12.280 33.830 12.700 34.040 ;
        RECT 13.170 33.830 13.590 34.040 ;
        RECT 14.400 33.870 15.860 34.040 ;
        RECT 12.350 33.770 12.610 33.830 ;
        RECT 13.260 33.770 13.520 33.830 ;
        RECT 14.860 33.810 15.150 33.870 ;
        RECT 16.380 33.700 16.800 34.040 ;
        RECT 17.060 34.000 17.230 34.870 ;
        RECT 17.610 34.000 17.780 34.690 ;
        RECT 21.750 34.650 21.920 35.340 ;
        RECT 22.290 34.480 22.460 35.350 ;
        RECT 22.730 35.310 23.150 35.590 ;
        RECT 24.370 35.480 24.540 35.810 ;
        RECT 25.990 35.520 26.250 35.610 ;
        RECT 26.900 35.520 27.160 35.610 ;
        RECT 23.670 35.310 25.090 35.480 ;
        RECT 25.900 35.310 26.320 35.520 ;
        RECT 26.830 35.310 27.250 35.520 ;
        RECT 22.730 34.870 24.310 35.040 ;
        RECT 25.520 34.920 25.690 35.250 ;
        RECT 19.560 34.100 19.730 34.430 ;
        RECT 20.970 34.310 22.550 34.480 ;
        RECT 18.030 33.830 18.450 34.040 ;
        RECT 18.920 33.830 19.340 34.040 ;
        RECT 20.150 33.870 21.610 34.040 ;
        RECT 18.100 33.770 18.360 33.830 ;
        RECT 19.010 33.770 19.270 33.830 ;
        RECT 20.610 33.810 20.900 33.870 ;
        RECT 22.130 33.700 22.550 34.040 ;
        RECT 22.810 34.000 22.980 34.870 ;
        RECT 23.360 34.000 23.530 34.690 ;
        RECT 27.500 34.650 27.670 35.340 ;
        RECT 28.040 34.480 28.210 35.350 ;
        RECT 28.480 35.310 28.900 35.590 ;
        RECT 30.120 35.480 30.290 35.810 ;
        RECT 31.740 35.520 32.000 35.610 ;
        RECT 32.650 35.520 32.910 35.610 ;
        RECT 29.420 35.310 30.840 35.480 ;
        RECT 31.650 35.310 32.070 35.520 ;
        RECT 32.580 35.310 33.000 35.520 ;
        RECT 28.480 34.870 30.060 35.040 ;
        RECT 31.270 34.920 31.440 35.250 ;
        RECT 25.310 34.100 25.480 34.430 ;
        RECT 26.720 34.310 28.300 34.480 ;
        RECT 23.780 33.830 24.200 34.040 ;
        RECT 24.670 33.830 25.090 34.040 ;
        RECT 25.900 33.870 27.360 34.040 ;
        RECT 23.850 33.770 24.110 33.830 ;
        RECT 24.760 33.770 25.020 33.830 ;
        RECT 26.360 33.810 26.650 33.870 ;
        RECT 27.880 33.700 28.300 34.040 ;
        RECT 28.560 34.000 28.730 34.870 ;
        RECT 29.110 34.000 29.280 34.690 ;
        RECT 33.250 34.650 33.420 35.340 ;
        RECT 33.790 34.480 33.960 35.350 ;
        RECT 34.230 35.310 34.650 35.590 ;
        RECT 35.870 35.480 36.040 35.810 ;
        RECT 37.490 35.520 37.750 35.610 ;
        RECT 38.400 35.520 38.660 35.610 ;
        RECT 35.170 35.310 36.590 35.480 ;
        RECT 37.400 35.310 37.820 35.520 ;
        RECT 38.330 35.310 38.750 35.520 ;
        RECT 34.230 34.870 35.810 35.040 ;
        RECT 37.020 34.920 37.190 35.250 ;
        RECT 31.060 34.100 31.230 34.430 ;
        RECT 32.470 34.310 34.050 34.480 ;
        RECT 29.530 33.830 29.950 34.040 ;
        RECT 30.420 33.830 30.840 34.040 ;
        RECT 31.650 33.870 33.110 34.040 ;
        RECT 29.600 33.770 29.860 33.830 ;
        RECT 30.510 33.770 30.770 33.830 ;
        RECT 32.110 33.810 32.400 33.870 ;
        RECT 33.630 33.700 34.050 34.040 ;
        RECT 34.310 34.000 34.480 34.870 ;
        RECT 34.860 34.000 35.030 34.690 ;
        RECT 39.000 34.650 39.170 35.340 ;
        RECT 39.540 34.480 39.710 35.350 ;
        RECT 39.980 35.310 40.400 35.590 ;
        RECT 41.620 35.480 41.790 35.810 ;
        RECT 43.240 35.520 43.500 35.610 ;
        RECT 44.150 35.520 44.410 35.610 ;
        RECT 40.920 35.310 42.340 35.480 ;
        RECT 43.150 35.310 43.570 35.520 ;
        RECT 44.080 35.310 44.500 35.520 ;
        RECT 39.980 34.870 41.560 35.040 ;
        RECT 42.770 34.920 42.940 35.250 ;
        RECT 36.810 34.100 36.980 34.430 ;
        RECT 38.220 34.310 39.800 34.480 ;
        RECT 35.280 33.830 35.700 34.040 ;
        RECT 36.170 33.830 36.590 34.040 ;
        RECT 37.400 33.870 38.860 34.040 ;
        RECT 35.350 33.770 35.610 33.830 ;
        RECT 36.260 33.770 36.520 33.830 ;
        RECT 37.860 33.810 38.150 33.870 ;
        RECT 39.380 33.700 39.800 34.040 ;
        RECT 40.060 34.000 40.230 34.870 ;
        RECT 40.610 34.000 40.780 34.690 ;
        RECT 44.750 34.650 44.920 35.340 ;
        RECT 45.290 34.480 45.460 35.350 ;
        RECT 45.730 35.310 46.150 35.590 ;
        RECT 47.370 35.480 47.540 35.810 ;
        RECT 48.990 35.520 49.250 35.610 ;
        RECT 49.900 35.520 50.160 35.610 ;
        RECT 46.670 35.310 48.090 35.480 ;
        RECT 48.900 35.310 49.320 35.520 ;
        RECT 49.830 35.310 50.250 35.520 ;
        RECT 45.730 34.870 47.310 35.040 ;
        RECT 48.520 34.920 48.690 35.250 ;
        RECT 42.560 34.100 42.730 34.430 ;
        RECT 43.970 34.310 45.550 34.480 ;
        RECT 41.030 33.830 41.450 34.040 ;
        RECT 41.920 33.830 42.340 34.040 ;
        RECT 43.150 33.870 44.610 34.040 ;
        RECT 41.100 33.770 41.360 33.830 ;
        RECT 42.010 33.770 42.270 33.830 ;
        RECT 43.610 33.810 43.900 33.870 ;
        RECT 45.130 33.700 45.550 34.040 ;
        RECT 45.810 34.000 45.980 34.870 ;
        RECT 46.360 34.000 46.530 34.690 ;
        RECT 50.500 34.650 50.670 35.340 ;
        RECT 51.040 34.480 51.210 35.350 ;
        RECT 51.480 35.310 51.900 35.590 ;
        RECT 53.120 35.480 53.290 35.810 ;
        RECT 54.740 35.520 55.000 35.610 ;
        RECT 55.650 35.520 55.910 35.610 ;
        RECT 52.420 35.310 53.840 35.480 ;
        RECT 54.650 35.310 55.070 35.520 ;
        RECT 55.580 35.310 56.000 35.520 ;
        RECT 51.480 34.870 53.060 35.040 ;
        RECT 54.270 34.920 54.440 35.250 ;
        RECT 48.310 34.100 48.480 34.430 ;
        RECT 49.720 34.310 51.300 34.480 ;
        RECT 46.780 33.830 47.200 34.040 ;
        RECT 47.670 33.830 48.090 34.040 ;
        RECT 48.900 33.870 50.360 34.040 ;
        RECT 46.850 33.770 47.110 33.830 ;
        RECT 47.760 33.770 48.020 33.830 ;
        RECT 49.360 33.810 49.650 33.870 ;
        RECT 50.880 33.700 51.300 34.040 ;
        RECT 51.560 34.000 51.730 34.870 ;
        RECT 52.110 34.000 52.280 34.690 ;
        RECT 56.250 34.650 56.420 35.340 ;
        RECT 56.790 34.480 56.960 35.350 ;
        RECT 57.230 35.310 57.650 35.590 ;
        RECT 58.870 35.480 59.040 35.810 ;
        RECT 60.490 35.520 60.750 35.610 ;
        RECT 61.400 35.520 61.660 35.610 ;
        RECT 58.170 35.310 59.590 35.480 ;
        RECT 60.400 35.310 60.820 35.520 ;
        RECT 61.330 35.310 61.750 35.520 ;
        RECT 57.230 34.870 58.810 35.040 ;
        RECT 60.020 34.920 60.190 35.250 ;
        RECT 54.060 34.100 54.230 34.430 ;
        RECT 55.470 34.310 57.050 34.480 ;
        RECT 52.530 33.830 52.950 34.040 ;
        RECT 53.420 33.830 53.840 34.040 ;
        RECT 54.650 33.870 56.110 34.040 ;
        RECT 52.600 33.770 52.860 33.830 ;
        RECT 53.510 33.770 53.770 33.830 ;
        RECT 55.110 33.810 55.400 33.870 ;
        RECT 56.630 33.700 57.050 34.040 ;
        RECT 57.310 34.000 57.480 34.870 ;
        RECT 57.860 34.000 58.030 34.690 ;
        RECT 62.000 34.650 62.170 35.340 ;
        RECT 62.540 34.480 62.710 35.350 ;
        RECT 62.980 35.310 63.400 35.590 ;
        RECT 64.620 35.480 64.790 35.810 ;
        RECT 66.240 35.520 66.500 35.610 ;
        RECT 67.150 35.520 67.410 35.610 ;
        RECT 63.920 35.310 65.340 35.480 ;
        RECT 66.150 35.310 66.570 35.520 ;
        RECT 67.080 35.310 67.500 35.520 ;
        RECT 62.980 34.870 64.560 35.040 ;
        RECT 65.770 34.920 65.940 35.250 ;
        RECT 59.810 34.100 59.980 34.430 ;
        RECT 61.220 34.310 62.800 34.480 ;
        RECT 58.280 33.830 58.700 34.040 ;
        RECT 59.170 33.830 59.590 34.040 ;
        RECT 60.400 33.870 61.860 34.040 ;
        RECT 58.350 33.770 58.610 33.830 ;
        RECT 59.260 33.770 59.520 33.830 ;
        RECT 60.860 33.810 61.150 33.870 ;
        RECT 62.380 33.700 62.800 34.040 ;
        RECT 63.060 34.000 63.230 34.870 ;
        RECT 63.610 34.000 63.780 34.690 ;
        RECT 67.750 34.650 67.920 35.340 ;
        RECT 68.290 34.480 68.460 35.350 ;
        RECT 68.730 35.310 69.150 35.590 ;
        RECT 70.370 35.480 70.540 35.810 ;
        RECT 71.990 35.520 72.250 35.610 ;
        RECT 72.900 35.520 73.160 35.610 ;
        RECT 69.670 35.310 71.090 35.480 ;
        RECT 71.900 35.310 72.320 35.520 ;
        RECT 72.830 35.310 73.250 35.520 ;
        RECT 68.730 34.870 70.310 35.040 ;
        RECT 71.520 34.920 71.690 35.250 ;
        RECT 65.560 34.100 65.730 34.430 ;
        RECT 66.970 34.310 68.550 34.480 ;
        RECT 64.030 33.830 64.450 34.040 ;
        RECT 64.920 33.830 65.340 34.040 ;
        RECT 66.150 33.870 67.610 34.040 ;
        RECT 64.100 33.770 64.360 33.830 ;
        RECT 65.010 33.770 65.270 33.830 ;
        RECT 66.610 33.810 66.900 33.870 ;
        RECT 68.130 33.700 68.550 34.040 ;
        RECT 68.810 34.000 68.980 34.870 ;
        RECT 69.360 34.000 69.530 34.690 ;
        RECT 73.500 34.650 73.670 35.340 ;
        RECT 74.040 34.480 74.210 35.350 ;
        RECT 74.480 35.310 74.900 35.590 ;
        RECT 76.120 35.480 76.290 35.810 ;
        RECT 77.740 35.520 78.000 35.610 ;
        RECT 78.650 35.520 78.910 35.610 ;
        RECT 75.420 35.310 76.840 35.480 ;
        RECT 77.650 35.310 78.070 35.520 ;
        RECT 78.580 35.310 79.000 35.520 ;
        RECT 74.480 34.870 76.060 35.040 ;
        RECT 77.270 34.920 77.440 35.250 ;
        RECT 71.310 34.100 71.480 34.430 ;
        RECT 72.720 34.310 74.300 34.480 ;
        RECT 69.780 33.830 70.200 34.040 ;
        RECT 70.670 33.830 71.090 34.040 ;
        RECT 71.900 33.870 73.360 34.040 ;
        RECT 69.850 33.770 70.110 33.830 ;
        RECT 70.760 33.770 71.020 33.830 ;
        RECT 72.360 33.810 72.650 33.870 ;
        RECT 73.880 33.700 74.300 34.040 ;
        RECT 74.560 34.000 74.730 34.870 ;
        RECT 75.110 34.000 75.280 34.690 ;
        RECT 79.250 34.650 79.420 35.340 ;
        RECT 79.790 34.480 79.960 35.350 ;
        RECT 80.230 35.310 80.650 35.590 ;
        RECT 81.870 35.480 82.040 35.810 ;
        RECT 83.490 35.520 83.750 35.610 ;
        RECT 84.400 35.520 84.660 35.610 ;
        RECT 81.170 35.310 82.590 35.480 ;
        RECT 83.400 35.310 83.820 35.520 ;
        RECT 84.330 35.310 84.750 35.520 ;
        RECT 80.230 34.870 81.810 35.040 ;
        RECT 83.020 34.920 83.190 35.250 ;
        RECT 77.060 34.100 77.230 34.430 ;
        RECT 78.470 34.310 80.050 34.480 ;
        RECT 75.530 33.830 75.950 34.040 ;
        RECT 76.420 33.830 76.840 34.040 ;
        RECT 77.650 33.870 79.110 34.040 ;
        RECT 75.600 33.770 75.860 33.830 ;
        RECT 76.510 33.770 76.770 33.830 ;
        RECT 78.110 33.810 78.400 33.870 ;
        RECT 79.630 33.700 80.050 34.040 ;
        RECT 80.310 34.000 80.480 34.870 ;
        RECT 80.860 34.000 81.030 34.690 ;
        RECT 85.000 34.650 85.170 35.340 ;
        RECT 85.540 34.480 85.710 35.350 ;
        RECT 85.980 35.310 86.400 35.590 ;
        RECT 87.620 35.480 87.790 35.810 ;
        RECT 89.240 35.520 89.500 35.610 ;
        RECT 90.150 35.520 90.410 35.610 ;
        RECT 86.920 35.310 88.340 35.480 ;
        RECT 89.150 35.310 89.570 35.520 ;
        RECT 90.080 35.310 90.500 35.520 ;
        RECT 85.980 34.870 87.560 35.040 ;
        RECT 88.770 34.920 88.940 35.250 ;
        RECT 82.810 34.100 82.980 34.430 ;
        RECT 84.220 34.310 85.800 34.480 ;
        RECT 81.280 33.830 81.700 34.040 ;
        RECT 82.170 33.830 82.590 34.040 ;
        RECT 83.400 33.870 84.860 34.040 ;
        RECT 81.350 33.770 81.610 33.830 ;
        RECT 82.260 33.770 82.520 33.830 ;
        RECT 83.860 33.810 84.150 33.870 ;
        RECT 85.380 33.700 85.800 34.040 ;
        RECT 86.060 34.000 86.230 34.870 ;
        RECT 86.610 34.000 86.780 34.690 ;
        RECT 90.750 34.650 90.920 35.340 ;
        RECT 91.290 34.480 91.460 35.350 ;
        RECT 91.730 35.310 92.150 35.590 ;
        RECT 93.370 35.480 93.540 35.810 ;
        RECT 92.670 35.310 94.090 35.480 ;
        RECT 91.730 34.870 93.310 35.040 ;
        RECT 88.560 34.100 88.730 34.430 ;
        RECT 89.970 34.310 91.550 34.480 ;
        RECT 87.030 33.830 87.450 34.040 ;
        RECT 87.920 33.830 88.340 34.040 ;
        RECT 89.150 33.870 90.610 34.040 ;
        RECT 87.100 33.770 87.360 33.830 ;
        RECT 88.010 33.770 88.270 33.830 ;
        RECT 89.610 33.810 89.900 33.870 ;
        RECT 91.130 33.700 91.550 34.040 ;
        RECT 91.810 34.000 91.980 34.870 ;
        RECT 92.360 34.000 92.530 34.690 ;
        RECT 94.310 34.100 94.480 34.430 ;
        RECT 92.780 33.830 93.200 34.040 ;
        RECT 93.670 33.830 94.090 34.040 ;
        RECT 92.850 33.770 93.110 33.830 ;
        RECT 93.760 33.770 94.020 33.830 ;
        RECT 2.990 33.110 3.250 33.200 ;
        RECT 3.900 33.110 4.160 33.200 ;
        RECT 2.900 32.900 3.320 33.110 ;
        RECT 3.830 32.900 4.250 33.110 ;
        RECT 2.520 32.510 2.690 32.840 ;
        RECT 4.500 32.240 4.670 32.930 ;
        RECT 5.040 32.070 5.210 32.940 ;
        RECT 5.480 32.900 5.900 33.180 ;
        RECT 7.120 33.070 7.290 33.400 ;
        RECT 8.740 33.110 9.000 33.200 ;
        RECT 9.650 33.110 9.910 33.200 ;
        RECT 6.420 32.900 7.840 33.070 ;
        RECT 8.650 32.900 9.070 33.110 ;
        RECT 9.580 32.900 10.000 33.110 ;
        RECT 5.480 32.460 7.060 32.630 ;
        RECT 8.270 32.510 8.440 32.840 ;
        RECT 3.720 31.900 5.300 32.070 ;
        RECT 2.900 31.460 4.360 31.630 ;
        RECT 3.360 31.400 3.650 31.460 ;
        RECT 4.880 31.290 5.300 31.630 ;
        RECT 5.560 31.590 5.730 32.460 ;
        RECT 6.110 31.590 6.280 32.280 ;
        RECT 10.250 32.240 10.420 32.930 ;
        RECT 10.790 32.070 10.960 32.940 ;
        RECT 11.230 32.900 11.650 33.180 ;
        RECT 12.870 33.070 13.040 33.400 ;
        RECT 14.490 33.110 14.750 33.200 ;
        RECT 15.400 33.110 15.660 33.200 ;
        RECT 12.170 32.900 13.590 33.070 ;
        RECT 14.400 32.900 14.820 33.110 ;
        RECT 15.330 32.900 15.750 33.110 ;
        RECT 11.230 32.460 12.810 32.630 ;
        RECT 14.020 32.510 14.190 32.840 ;
        RECT 8.060 31.690 8.230 32.020 ;
        RECT 9.470 31.900 11.050 32.070 ;
        RECT 6.530 31.420 6.950 31.630 ;
        RECT 7.420 31.420 7.840 31.630 ;
        RECT 8.650 31.460 10.110 31.630 ;
        RECT 6.600 31.360 6.860 31.420 ;
        RECT 7.510 31.360 7.770 31.420 ;
        RECT 9.110 31.400 9.400 31.460 ;
        RECT 10.630 31.290 11.050 31.630 ;
        RECT 11.310 31.590 11.480 32.460 ;
        RECT 11.860 31.590 12.030 32.280 ;
        RECT 16.000 32.240 16.170 32.930 ;
        RECT 16.540 32.070 16.710 32.940 ;
        RECT 16.980 32.900 17.400 33.180 ;
        RECT 18.620 33.070 18.790 33.400 ;
        RECT 20.240 33.110 20.500 33.200 ;
        RECT 21.150 33.110 21.410 33.200 ;
        RECT 17.920 32.900 19.340 33.070 ;
        RECT 20.150 32.900 20.570 33.110 ;
        RECT 21.080 32.900 21.500 33.110 ;
        RECT 16.980 32.460 18.560 32.630 ;
        RECT 19.770 32.510 19.940 32.840 ;
        RECT 13.810 31.690 13.980 32.020 ;
        RECT 15.220 31.900 16.800 32.070 ;
        RECT 12.280 31.420 12.700 31.630 ;
        RECT 13.170 31.420 13.590 31.630 ;
        RECT 14.400 31.460 15.860 31.630 ;
        RECT 12.350 31.360 12.610 31.420 ;
        RECT 13.260 31.360 13.520 31.420 ;
        RECT 14.860 31.400 15.150 31.460 ;
        RECT 16.380 31.290 16.800 31.630 ;
        RECT 17.060 31.590 17.230 32.460 ;
        RECT 17.610 31.590 17.780 32.280 ;
        RECT 21.750 32.240 21.920 32.930 ;
        RECT 22.290 32.070 22.460 32.940 ;
        RECT 22.730 32.900 23.150 33.180 ;
        RECT 24.370 33.070 24.540 33.400 ;
        RECT 25.990 33.110 26.250 33.200 ;
        RECT 26.900 33.110 27.160 33.200 ;
        RECT 23.670 32.900 25.090 33.070 ;
        RECT 25.900 32.900 26.320 33.110 ;
        RECT 26.830 32.900 27.250 33.110 ;
        RECT 22.730 32.460 24.310 32.630 ;
        RECT 25.520 32.510 25.690 32.840 ;
        RECT 19.560 31.690 19.730 32.020 ;
        RECT 20.970 31.900 22.550 32.070 ;
        RECT 18.030 31.420 18.450 31.630 ;
        RECT 18.920 31.420 19.340 31.630 ;
        RECT 20.150 31.460 21.610 31.630 ;
        RECT 18.100 31.360 18.360 31.420 ;
        RECT 19.010 31.360 19.270 31.420 ;
        RECT 20.610 31.400 20.900 31.460 ;
        RECT 22.130 31.290 22.550 31.630 ;
        RECT 22.810 31.590 22.980 32.460 ;
        RECT 23.360 31.590 23.530 32.280 ;
        RECT 27.500 32.240 27.670 32.930 ;
        RECT 28.040 32.070 28.210 32.940 ;
        RECT 28.480 32.900 28.900 33.180 ;
        RECT 30.120 33.070 30.290 33.400 ;
        RECT 31.740 33.110 32.000 33.200 ;
        RECT 32.650 33.110 32.910 33.200 ;
        RECT 29.420 32.900 30.840 33.070 ;
        RECT 31.650 32.900 32.070 33.110 ;
        RECT 32.580 32.900 33.000 33.110 ;
        RECT 28.480 32.460 30.060 32.630 ;
        RECT 31.270 32.510 31.440 32.840 ;
        RECT 25.310 31.690 25.480 32.020 ;
        RECT 26.720 31.900 28.300 32.070 ;
        RECT 23.780 31.420 24.200 31.630 ;
        RECT 24.670 31.420 25.090 31.630 ;
        RECT 25.900 31.460 27.360 31.630 ;
        RECT 23.850 31.360 24.110 31.420 ;
        RECT 24.760 31.360 25.020 31.420 ;
        RECT 26.360 31.400 26.650 31.460 ;
        RECT 27.880 31.290 28.300 31.630 ;
        RECT 28.560 31.590 28.730 32.460 ;
        RECT 29.110 31.590 29.280 32.280 ;
        RECT 33.250 32.240 33.420 32.930 ;
        RECT 33.790 32.070 33.960 32.940 ;
        RECT 34.230 32.900 34.650 33.180 ;
        RECT 35.870 33.070 36.040 33.400 ;
        RECT 37.490 33.110 37.750 33.200 ;
        RECT 38.400 33.110 38.660 33.200 ;
        RECT 35.170 32.900 36.590 33.070 ;
        RECT 37.400 32.900 37.820 33.110 ;
        RECT 38.330 32.900 38.750 33.110 ;
        RECT 34.230 32.460 35.810 32.630 ;
        RECT 37.020 32.510 37.190 32.840 ;
        RECT 31.060 31.690 31.230 32.020 ;
        RECT 32.470 31.900 34.050 32.070 ;
        RECT 29.530 31.420 29.950 31.630 ;
        RECT 30.420 31.420 30.840 31.630 ;
        RECT 31.650 31.460 33.110 31.630 ;
        RECT 29.600 31.360 29.860 31.420 ;
        RECT 30.510 31.360 30.770 31.420 ;
        RECT 32.110 31.400 32.400 31.460 ;
        RECT 33.630 31.290 34.050 31.630 ;
        RECT 34.310 31.590 34.480 32.460 ;
        RECT 34.860 31.590 35.030 32.280 ;
        RECT 39.000 32.240 39.170 32.930 ;
        RECT 39.540 32.070 39.710 32.940 ;
        RECT 39.980 32.900 40.400 33.180 ;
        RECT 41.620 33.070 41.790 33.400 ;
        RECT 43.240 33.110 43.500 33.200 ;
        RECT 44.150 33.110 44.410 33.200 ;
        RECT 40.920 32.900 42.340 33.070 ;
        RECT 43.150 32.900 43.570 33.110 ;
        RECT 44.080 32.900 44.500 33.110 ;
        RECT 39.980 32.460 41.560 32.630 ;
        RECT 42.770 32.510 42.940 32.840 ;
        RECT 36.810 31.690 36.980 32.020 ;
        RECT 38.220 31.900 39.800 32.070 ;
        RECT 35.280 31.420 35.700 31.630 ;
        RECT 36.170 31.420 36.590 31.630 ;
        RECT 37.400 31.460 38.860 31.630 ;
        RECT 35.350 31.360 35.610 31.420 ;
        RECT 36.260 31.360 36.520 31.420 ;
        RECT 37.860 31.400 38.150 31.460 ;
        RECT 39.380 31.290 39.800 31.630 ;
        RECT 40.060 31.590 40.230 32.460 ;
        RECT 40.610 31.590 40.780 32.280 ;
        RECT 44.750 32.240 44.920 32.930 ;
        RECT 45.290 32.070 45.460 32.940 ;
        RECT 45.730 32.900 46.150 33.180 ;
        RECT 47.370 33.070 47.540 33.400 ;
        RECT 48.990 33.110 49.250 33.200 ;
        RECT 49.900 33.110 50.160 33.200 ;
        RECT 46.670 32.900 48.090 33.070 ;
        RECT 48.900 32.900 49.320 33.110 ;
        RECT 49.830 32.900 50.250 33.110 ;
        RECT 45.730 32.460 47.310 32.630 ;
        RECT 48.520 32.510 48.690 32.840 ;
        RECT 42.560 31.690 42.730 32.020 ;
        RECT 43.970 31.900 45.550 32.070 ;
        RECT 41.030 31.420 41.450 31.630 ;
        RECT 41.920 31.420 42.340 31.630 ;
        RECT 43.150 31.460 44.610 31.630 ;
        RECT 41.100 31.360 41.360 31.420 ;
        RECT 42.010 31.360 42.270 31.420 ;
        RECT 43.610 31.400 43.900 31.460 ;
        RECT 45.130 31.290 45.550 31.630 ;
        RECT 45.810 31.590 45.980 32.460 ;
        RECT 46.360 31.590 46.530 32.280 ;
        RECT 50.500 32.240 50.670 32.930 ;
        RECT 51.040 32.070 51.210 32.940 ;
        RECT 51.480 32.900 51.900 33.180 ;
        RECT 53.120 33.070 53.290 33.400 ;
        RECT 54.740 33.110 55.000 33.200 ;
        RECT 55.650 33.110 55.910 33.200 ;
        RECT 52.420 32.900 53.840 33.070 ;
        RECT 54.650 32.900 55.070 33.110 ;
        RECT 55.580 32.900 56.000 33.110 ;
        RECT 51.480 32.460 53.060 32.630 ;
        RECT 54.270 32.510 54.440 32.840 ;
        RECT 48.310 31.690 48.480 32.020 ;
        RECT 49.720 31.900 51.300 32.070 ;
        RECT 46.780 31.420 47.200 31.630 ;
        RECT 47.670 31.420 48.090 31.630 ;
        RECT 48.900 31.460 50.360 31.630 ;
        RECT 46.850 31.360 47.110 31.420 ;
        RECT 47.760 31.360 48.020 31.420 ;
        RECT 49.360 31.400 49.650 31.460 ;
        RECT 50.880 31.290 51.300 31.630 ;
        RECT 51.560 31.590 51.730 32.460 ;
        RECT 52.110 31.590 52.280 32.280 ;
        RECT 56.250 32.240 56.420 32.930 ;
        RECT 56.790 32.070 56.960 32.940 ;
        RECT 57.230 32.900 57.650 33.180 ;
        RECT 58.870 33.070 59.040 33.400 ;
        RECT 60.490 33.110 60.750 33.200 ;
        RECT 61.400 33.110 61.660 33.200 ;
        RECT 58.170 32.900 59.590 33.070 ;
        RECT 60.400 32.900 60.820 33.110 ;
        RECT 61.330 32.900 61.750 33.110 ;
        RECT 57.230 32.460 58.810 32.630 ;
        RECT 60.020 32.510 60.190 32.840 ;
        RECT 54.060 31.690 54.230 32.020 ;
        RECT 55.470 31.900 57.050 32.070 ;
        RECT 52.530 31.420 52.950 31.630 ;
        RECT 53.420 31.420 53.840 31.630 ;
        RECT 54.650 31.460 56.110 31.630 ;
        RECT 52.600 31.360 52.860 31.420 ;
        RECT 53.510 31.360 53.770 31.420 ;
        RECT 55.110 31.400 55.400 31.460 ;
        RECT 56.630 31.290 57.050 31.630 ;
        RECT 57.310 31.590 57.480 32.460 ;
        RECT 57.860 31.590 58.030 32.280 ;
        RECT 62.000 32.240 62.170 32.930 ;
        RECT 62.540 32.070 62.710 32.940 ;
        RECT 62.980 32.900 63.400 33.180 ;
        RECT 64.620 33.070 64.790 33.400 ;
        RECT 66.240 33.110 66.500 33.200 ;
        RECT 67.150 33.110 67.410 33.200 ;
        RECT 63.920 32.900 65.340 33.070 ;
        RECT 66.150 32.900 66.570 33.110 ;
        RECT 67.080 32.900 67.500 33.110 ;
        RECT 62.980 32.460 64.560 32.630 ;
        RECT 65.770 32.510 65.940 32.840 ;
        RECT 59.810 31.690 59.980 32.020 ;
        RECT 61.220 31.900 62.800 32.070 ;
        RECT 58.280 31.420 58.700 31.630 ;
        RECT 59.170 31.420 59.590 31.630 ;
        RECT 60.400 31.460 61.860 31.630 ;
        RECT 58.350 31.360 58.610 31.420 ;
        RECT 59.260 31.360 59.520 31.420 ;
        RECT 60.860 31.400 61.150 31.460 ;
        RECT 62.380 31.290 62.800 31.630 ;
        RECT 63.060 31.590 63.230 32.460 ;
        RECT 63.610 31.590 63.780 32.280 ;
        RECT 67.750 32.240 67.920 32.930 ;
        RECT 68.290 32.070 68.460 32.940 ;
        RECT 68.730 32.900 69.150 33.180 ;
        RECT 70.370 33.070 70.540 33.400 ;
        RECT 71.990 33.110 72.250 33.200 ;
        RECT 72.900 33.110 73.160 33.200 ;
        RECT 69.670 32.900 71.090 33.070 ;
        RECT 71.900 32.900 72.320 33.110 ;
        RECT 72.830 32.900 73.250 33.110 ;
        RECT 68.730 32.460 70.310 32.630 ;
        RECT 71.520 32.510 71.690 32.840 ;
        RECT 65.560 31.690 65.730 32.020 ;
        RECT 66.970 31.900 68.550 32.070 ;
        RECT 64.030 31.420 64.450 31.630 ;
        RECT 64.920 31.420 65.340 31.630 ;
        RECT 66.150 31.460 67.610 31.630 ;
        RECT 64.100 31.360 64.360 31.420 ;
        RECT 65.010 31.360 65.270 31.420 ;
        RECT 66.610 31.400 66.900 31.460 ;
        RECT 68.130 31.290 68.550 31.630 ;
        RECT 68.810 31.590 68.980 32.460 ;
        RECT 69.360 31.590 69.530 32.280 ;
        RECT 73.500 32.240 73.670 32.930 ;
        RECT 74.040 32.070 74.210 32.940 ;
        RECT 74.480 32.900 74.900 33.180 ;
        RECT 76.120 33.070 76.290 33.400 ;
        RECT 77.740 33.110 78.000 33.200 ;
        RECT 78.650 33.110 78.910 33.200 ;
        RECT 75.420 32.900 76.840 33.070 ;
        RECT 77.650 32.900 78.070 33.110 ;
        RECT 78.580 32.900 79.000 33.110 ;
        RECT 74.480 32.460 76.060 32.630 ;
        RECT 77.270 32.510 77.440 32.840 ;
        RECT 71.310 31.690 71.480 32.020 ;
        RECT 72.720 31.900 74.300 32.070 ;
        RECT 69.780 31.420 70.200 31.630 ;
        RECT 70.670 31.420 71.090 31.630 ;
        RECT 71.900 31.460 73.360 31.630 ;
        RECT 69.850 31.360 70.110 31.420 ;
        RECT 70.760 31.360 71.020 31.420 ;
        RECT 72.360 31.400 72.650 31.460 ;
        RECT 73.880 31.290 74.300 31.630 ;
        RECT 74.560 31.590 74.730 32.460 ;
        RECT 75.110 31.590 75.280 32.280 ;
        RECT 79.250 32.240 79.420 32.930 ;
        RECT 79.790 32.070 79.960 32.940 ;
        RECT 80.230 32.900 80.650 33.180 ;
        RECT 81.870 33.070 82.040 33.400 ;
        RECT 83.490 33.110 83.750 33.200 ;
        RECT 84.400 33.110 84.660 33.200 ;
        RECT 81.170 32.900 82.590 33.070 ;
        RECT 83.400 32.900 83.820 33.110 ;
        RECT 84.330 32.900 84.750 33.110 ;
        RECT 80.230 32.460 81.810 32.630 ;
        RECT 83.020 32.510 83.190 32.840 ;
        RECT 77.060 31.690 77.230 32.020 ;
        RECT 78.470 31.900 80.050 32.070 ;
        RECT 75.530 31.420 75.950 31.630 ;
        RECT 76.420 31.420 76.840 31.630 ;
        RECT 77.650 31.460 79.110 31.630 ;
        RECT 75.600 31.360 75.860 31.420 ;
        RECT 76.510 31.360 76.770 31.420 ;
        RECT 78.110 31.400 78.400 31.460 ;
        RECT 79.630 31.290 80.050 31.630 ;
        RECT 80.310 31.590 80.480 32.460 ;
        RECT 80.860 31.590 81.030 32.280 ;
        RECT 85.000 32.240 85.170 32.930 ;
        RECT 85.540 32.070 85.710 32.940 ;
        RECT 85.980 32.900 86.400 33.180 ;
        RECT 87.620 33.070 87.790 33.400 ;
        RECT 89.240 33.110 89.500 33.200 ;
        RECT 90.150 33.110 90.410 33.200 ;
        RECT 86.920 32.900 88.340 33.070 ;
        RECT 89.150 32.900 89.570 33.110 ;
        RECT 90.080 32.900 90.500 33.110 ;
        RECT 85.980 32.460 87.560 32.630 ;
        RECT 88.770 32.510 88.940 32.840 ;
        RECT 82.810 31.690 82.980 32.020 ;
        RECT 84.220 31.900 85.800 32.070 ;
        RECT 81.280 31.420 81.700 31.630 ;
        RECT 82.170 31.420 82.590 31.630 ;
        RECT 83.400 31.460 84.860 31.630 ;
        RECT 81.350 31.360 81.610 31.420 ;
        RECT 82.260 31.360 82.520 31.420 ;
        RECT 83.860 31.400 84.150 31.460 ;
        RECT 85.380 31.290 85.800 31.630 ;
        RECT 86.060 31.590 86.230 32.460 ;
        RECT 86.610 31.590 86.780 32.280 ;
        RECT 90.750 32.240 90.920 32.930 ;
        RECT 91.290 32.070 91.460 32.940 ;
        RECT 91.730 32.900 92.150 33.180 ;
        RECT 93.370 33.070 93.540 33.400 ;
        RECT 92.670 32.900 94.090 33.070 ;
        RECT 91.730 32.460 93.310 32.630 ;
        RECT 88.560 31.690 88.730 32.020 ;
        RECT 89.970 31.900 91.550 32.070 ;
        RECT 87.030 31.420 87.450 31.630 ;
        RECT 87.920 31.420 88.340 31.630 ;
        RECT 89.150 31.460 90.610 31.630 ;
        RECT 87.100 31.360 87.360 31.420 ;
        RECT 88.010 31.360 88.270 31.420 ;
        RECT 89.610 31.400 89.900 31.460 ;
        RECT 91.130 31.290 91.550 31.630 ;
        RECT 91.810 31.590 91.980 32.460 ;
        RECT 92.360 31.590 92.530 32.280 ;
        RECT 94.310 31.690 94.480 32.020 ;
        RECT 92.780 31.420 93.200 31.630 ;
        RECT 93.670 31.420 94.090 31.630 ;
        RECT 92.850 31.360 93.110 31.420 ;
        RECT 93.760 31.360 94.020 31.420 ;
        RECT 2.990 30.700 3.250 30.790 ;
        RECT 3.900 30.700 4.160 30.790 ;
        RECT 2.900 30.490 3.320 30.700 ;
        RECT 3.830 30.490 4.250 30.700 ;
        RECT 2.520 30.100 2.690 30.430 ;
        RECT 4.500 29.830 4.670 30.520 ;
        RECT 5.040 29.660 5.210 30.530 ;
        RECT 5.480 30.490 5.900 30.770 ;
        RECT 7.120 30.660 7.290 30.990 ;
        RECT 8.740 30.700 9.000 30.790 ;
        RECT 9.650 30.700 9.910 30.790 ;
        RECT 6.420 30.490 7.840 30.660 ;
        RECT 8.650 30.490 9.070 30.700 ;
        RECT 9.580 30.490 10.000 30.700 ;
        RECT 5.480 30.050 7.060 30.220 ;
        RECT 8.270 30.100 8.440 30.430 ;
        RECT 3.720 29.490 5.300 29.660 ;
        RECT 2.900 29.050 4.360 29.220 ;
        RECT 3.020 28.170 3.190 29.050 ;
        RECT 3.360 28.990 3.650 29.050 ;
        RECT 4.880 28.880 5.300 29.220 ;
        RECT 5.560 29.180 5.730 30.050 ;
        RECT 6.110 29.180 6.280 29.870 ;
        RECT 10.250 29.830 10.420 30.520 ;
        RECT 10.790 29.660 10.960 30.530 ;
        RECT 11.230 30.490 11.650 30.770 ;
        RECT 12.870 30.660 13.040 30.990 ;
        RECT 14.490 30.700 14.750 30.790 ;
        RECT 15.400 30.700 15.660 30.790 ;
        RECT 12.170 30.490 13.590 30.660 ;
        RECT 14.400 30.490 14.820 30.700 ;
        RECT 15.330 30.490 15.750 30.700 ;
        RECT 11.230 30.050 12.810 30.220 ;
        RECT 14.020 30.100 14.190 30.430 ;
        RECT 8.060 29.280 8.230 29.610 ;
        RECT 9.470 29.490 11.050 29.660 ;
        RECT 6.530 29.010 6.950 29.220 ;
        RECT 7.420 29.010 7.840 29.220 ;
        RECT 8.650 29.050 10.110 29.220 ;
        RECT 6.600 28.950 6.860 29.010 ;
        RECT 7.510 28.950 7.770 29.010 ;
        RECT 5.010 28.170 5.180 28.880 ;
        RECT 2.990 27.890 3.250 27.980 ;
        RECT 3.900 27.890 4.160 27.980 ;
        RECT 2.900 27.680 3.320 27.890 ;
        RECT 3.830 27.680 4.250 27.890 ;
        RECT 2.520 27.290 2.690 27.620 ;
        RECT 4.500 27.020 4.670 27.710 ;
        RECT 5.040 26.850 5.210 27.720 ;
        RECT 5.480 27.680 5.900 27.960 ;
        RECT 7.120 27.850 7.290 28.260 ;
        RECT 8.770 28.170 8.940 29.050 ;
        RECT 9.110 28.990 9.400 29.050 ;
        RECT 10.630 28.880 11.050 29.220 ;
        RECT 11.310 29.180 11.480 30.050 ;
        RECT 11.860 29.180 12.030 29.870 ;
        RECT 16.000 29.830 16.170 30.520 ;
        RECT 16.540 29.660 16.710 30.530 ;
        RECT 16.980 30.490 17.400 30.770 ;
        RECT 18.620 30.660 18.790 30.990 ;
        RECT 20.240 30.700 20.500 30.790 ;
        RECT 21.150 30.700 21.410 30.790 ;
        RECT 17.920 30.490 19.340 30.660 ;
        RECT 20.150 30.490 20.570 30.700 ;
        RECT 21.080 30.490 21.500 30.700 ;
        RECT 16.980 30.050 18.560 30.220 ;
        RECT 19.770 30.100 19.940 30.430 ;
        RECT 13.810 29.280 13.980 29.610 ;
        RECT 15.220 29.490 16.800 29.660 ;
        RECT 12.280 29.010 12.700 29.220 ;
        RECT 13.170 29.010 13.590 29.220 ;
        RECT 14.400 29.050 15.860 29.220 ;
        RECT 12.350 28.950 12.610 29.010 ;
        RECT 13.260 28.950 13.520 29.010 ;
        RECT 10.770 28.170 10.940 28.880 ;
        RECT 8.740 27.890 9.000 27.980 ;
        RECT 9.650 27.890 9.910 27.980 ;
        RECT 6.420 27.680 7.840 27.850 ;
        RECT 8.650 27.680 9.070 27.890 ;
        RECT 9.580 27.680 10.000 27.890 ;
        RECT 5.480 27.240 7.060 27.410 ;
        RECT 8.270 27.290 8.440 27.620 ;
        RECT 3.720 26.680 5.300 26.850 ;
        RECT 2.900 26.240 4.360 26.410 ;
        RECT 3.360 26.180 3.650 26.240 ;
        RECT 4.880 26.070 5.300 26.410 ;
        RECT 5.560 26.370 5.730 27.240 ;
        RECT 6.110 26.370 6.280 27.060 ;
        RECT 10.250 27.020 10.420 27.710 ;
        RECT 10.790 26.850 10.960 27.720 ;
        RECT 11.230 27.680 11.650 27.960 ;
        RECT 12.870 27.850 13.040 28.260 ;
        RECT 14.520 28.170 14.690 29.050 ;
        RECT 14.860 28.990 15.150 29.050 ;
        RECT 16.380 28.880 16.800 29.220 ;
        RECT 17.060 29.180 17.230 30.050 ;
        RECT 17.610 29.180 17.780 29.870 ;
        RECT 21.750 29.830 21.920 30.520 ;
        RECT 22.290 29.660 22.460 30.530 ;
        RECT 22.730 30.490 23.150 30.770 ;
        RECT 24.370 30.660 24.540 30.990 ;
        RECT 25.990 30.700 26.250 30.790 ;
        RECT 26.900 30.700 27.160 30.790 ;
        RECT 23.670 30.490 25.090 30.660 ;
        RECT 25.900 30.490 26.320 30.700 ;
        RECT 26.830 30.490 27.250 30.700 ;
        RECT 22.730 30.050 24.310 30.220 ;
        RECT 25.520 30.100 25.690 30.430 ;
        RECT 19.560 29.280 19.730 29.610 ;
        RECT 20.970 29.490 22.550 29.660 ;
        RECT 18.030 29.010 18.450 29.220 ;
        RECT 18.920 29.010 19.340 29.220 ;
        RECT 20.150 29.050 21.610 29.220 ;
        RECT 18.100 28.950 18.360 29.010 ;
        RECT 19.010 28.950 19.270 29.010 ;
        RECT 16.520 28.170 16.690 28.880 ;
        RECT 14.490 27.890 14.750 27.980 ;
        RECT 15.400 27.890 15.660 27.980 ;
        RECT 12.170 27.680 13.590 27.850 ;
        RECT 14.400 27.680 14.820 27.890 ;
        RECT 15.330 27.680 15.750 27.890 ;
        RECT 11.230 27.240 12.810 27.410 ;
        RECT 14.020 27.290 14.190 27.620 ;
        RECT 8.060 26.470 8.230 26.800 ;
        RECT 9.470 26.680 11.050 26.850 ;
        RECT 6.530 26.200 6.950 26.410 ;
        RECT 7.420 26.200 7.840 26.410 ;
        RECT 8.650 26.240 10.110 26.410 ;
        RECT 6.600 26.140 6.860 26.200 ;
        RECT 7.510 26.140 7.770 26.200 ;
        RECT 9.110 26.180 9.400 26.240 ;
        RECT 10.630 26.070 11.050 26.410 ;
        RECT 11.310 26.370 11.480 27.240 ;
        RECT 11.860 26.370 12.030 27.060 ;
        RECT 16.000 27.020 16.170 27.710 ;
        RECT 16.540 26.850 16.710 27.720 ;
        RECT 16.980 27.680 17.400 27.960 ;
        RECT 18.620 27.850 18.790 28.260 ;
        RECT 20.270 28.170 20.440 29.050 ;
        RECT 20.610 28.990 20.900 29.050 ;
        RECT 22.130 28.880 22.550 29.220 ;
        RECT 22.810 29.180 22.980 30.050 ;
        RECT 23.360 29.180 23.530 29.870 ;
        RECT 27.500 29.830 27.670 30.520 ;
        RECT 28.040 29.660 28.210 30.530 ;
        RECT 28.480 30.490 28.900 30.770 ;
        RECT 30.120 30.660 30.290 30.990 ;
        RECT 31.740 30.700 32.000 30.790 ;
        RECT 32.650 30.700 32.910 30.790 ;
        RECT 29.420 30.490 30.840 30.660 ;
        RECT 31.650 30.490 32.070 30.700 ;
        RECT 32.580 30.490 33.000 30.700 ;
        RECT 28.480 30.050 30.060 30.220 ;
        RECT 31.270 30.100 31.440 30.430 ;
        RECT 25.310 29.280 25.480 29.610 ;
        RECT 26.720 29.490 28.300 29.660 ;
        RECT 23.780 29.010 24.200 29.220 ;
        RECT 24.670 29.010 25.090 29.220 ;
        RECT 25.900 29.050 27.360 29.220 ;
        RECT 23.850 28.950 24.110 29.010 ;
        RECT 24.760 28.950 25.020 29.010 ;
        RECT 22.270 28.170 22.440 28.880 ;
        RECT 20.240 27.890 20.500 27.980 ;
        RECT 21.150 27.890 21.410 27.980 ;
        RECT 17.920 27.680 19.340 27.850 ;
        RECT 20.150 27.680 20.570 27.890 ;
        RECT 21.080 27.680 21.500 27.890 ;
        RECT 16.980 27.240 18.560 27.410 ;
        RECT 19.770 27.290 19.940 27.620 ;
        RECT 13.810 26.470 13.980 26.800 ;
        RECT 15.220 26.680 16.800 26.850 ;
        RECT 12.280 26.200 12.700 26.410 ;
        RECT 13.170 26.200 13.590 26.410 ;
        RECT 14.400 26.240 15.860 26.410 ;
        RECT 12.350 26.140 12.610 26.200 ;
        RECT 13.260 26.140 13.520 26.200 ;
        RECT 14.860 26.180 15.150 26.240 ;
        RECT 16.380 26.070 16.800 26.410 ;
        RECT 17.060 26.370 17.230 27.240 ;
        RECT 17.610 26.370 17.780 27.060 ;
        RECT 21.750 27.020 21.920 27.710 ;
        RECT 22.290 26.850 22.460 27.720 ;
        RECT 22.730 27.680 23.150 27.960 ;
        RECT 24.370 27.850 24.540 28.260 ;
        RECT 26.020 28.170 26.190 29.050 ;
        RECT 26.360 28.990 26.650 29.050 ;
        RECT 27.880 28.880 28.300 29.220 ;
        RECT 28.560 29.180 28.730 30.050 ;
        RECT 29.110 29.180 29.280 29.870 ;
        RECT 33.250 29.830 33.420 30.520 ;
        RECT 33.790 29.660 33.960 30.530 ;
        RECT 34.230 30.490 34.650 30.770 ;
        RECT 35.870 30.660 36.040 30.990 ;
        RECT 37.490 30.700 37.750 30.790 ;
        RECT 38.400 30.700 38.660 30.790 ;
        RECT 35.170 30.490 36.590 30.660 ;
        RECT 37.400 30.490 37.820 30.700 ;
        RECT 38.330 30.490 38.750 30.700 ;
        RECT 34.230 30.050 35.810 30.220 ;
        RECT 37.020 30.100 37.190 30.430 ;
        RECT 31.060 29.280 31.230 29.610 ;
        RECT 32.470 29.490 34.050 29.660 ;
        RECT 29.530 29.010 29.950 29.220 ;
        RECT 30.420 29.010 30.840 29.220 ;
        RECT 31.650 29.050 33.110 29.220 ;
        RECT 29.600 28.950 29.860 29.010 ;
        RECT 30.510 28.950 30.770 29.010 ;
        RECT 28.020 28.170 28.190 28.880 ;
        RECT 25.990 27.890 26.250 27.980 ;
        RECT 26.900 27.890 27.160 27.980 ;
        RECT 23.670 27.680 25.090 27.850 ;
        RECT 25.900 27.680 26.320 27.890 ;
        RECT 26.830 27.680 27.250 27.890 ;
        RECT 22.730 27.240 24.310 27.410 ;
        RECT 25.520 27.290 25.690 27.620 ;
        RECT 19.560 26.470 19.730 26.800 ;
        RECT 20.970 26.680 22.550 26.850 ;
        RECT 18.030 26.200 18.450 26.410 ;
        RECT 18.920 26.200 19.340 26.410 ;
        RECT 20.150 26.240 21.610 26.410 ;
        RECT 18.100 26.140 18.360 26.200 ;
        RECT 19.010 26.140 19.270 26.200 ;
        RECT 20.610 26.180 20.900 26.240 ;
        RECT 22.130 26.070 22.550 26.410 ;
        RECT 22.810 26.370 22.980 27.240 ;
        RECT 23.360 26.370 23.530 27.060 ;
        RECT 27.500 27.020 27.670 27.710 ;
        RECT 28.040 26.850 28.210 27.720 ;
        RECT 28.480 27.680 28.900 27.960 ;
        RECT 30.120 27.850 30.290 28.260 ;
        RECT 31.770 28.170 31.940 29.050 ;
        RECT 32.110 28.990 32.400 29.050 ;
        RECT 33.630 28.880 34.050 29.220 ;
        RECT 34.310 29.180 34.480 30.050 ;
        RECT 34.860 29.180 35.030 29.870 ;
        RECT 39.000 29.830 39.170 30.520 ;
        RECT 39.540 29.660 39.710 30.530 ;
        RECT 39.980 30.490 40.400 30.770 ;
        RECT 41.620 30.660 41.790 30.990 ;
        RECT 43.240 30.700 43.500 30.790 ;
        RECT 44.150 30.700 44.410 30.790 ;
        RECT 40.920 30.490 42.340 30.660 ;
        RECT 43.150 30.490 43.570 30.700 ;
        RECT 44.080 30.490 44.500 30.700 ;
        RECT 39.980 30.050 41.560 30.220 ;
        RECT 42.770 30.100 42.940 30.430 ;
        RECT 36.810 29.280 36.980 29.610 ;
        RECT 38.220 29.490 39.800 29.660 ;
        RECT 35.280 29.010 35.700 29.220 ;
        RECT 36.170 29.010 36.590 29.220 ;
        RECT 37.400 29.050 38.860 29.220 ;
        RECT 35.350 28.950 35.610 29.010 ;
        RECT 36.260 28.950 36.520 29.010 ;
        RECT 33.770 28.170 33.940 28.880 ;
        RECT 31.740 27.890 32.000 27.980 ;
        RECT 32.650 27.890 32.910 27.980 ;
        RECT 29.420 27.680 30.840 27.850 ;
        RECT 31.650 27.680 32.070 27.890 ;
        RECT 32.580 27.680 33.000 27.890 ;
        RECT 28.480 27.240 30.060 27.410 ;
        RECT 31.270 27.290 31.440 27.620 ;
        RECT 25.310 26.470 25.480 26.800 ;
        RECT 26.720 26.680 28.300 26.850 ;
        RECT 23.780 26.200 24.200 26.410 ;
        RECT 24.670 26.200 25.090 26.410 ;
        RECT 25.900 26.240 27.360 26.410 ;
        RECT 23.850 26.140 24.110 26.200 ;
        RECT 24.760 26.140 25.020 26.200 ;
        RECT 26.360 26.180 26.650 26.240 ;
        RECT 27.880 26.070 28.300 26.410 ;
        RECT 28.560 26.370 28.730 27.240 ;
        RECT 29.110 26.370 29.280 27.060 ;
        RECT 33.250 27.020 33.420 27.710 ;
        RECT 33.790 26.850 33.960 27.720 ;
        RECT 34.230 27.680 34.650 27.960 ;
        RECT 35.870 27.850 36.040 28.260 ;
        RECT 37.520 28.170 37.690 29.050 ;
        RECT 37.860 28.990 38.150 29.050 ;
        RECT 39.380 28.880 39.800 29.220 ;
        RECT 40.060 29.180 40.230 30.050 ;
        RECT 40.610 29.180 40.780 29.870 ;
        RECT 44.750 29.830 44.920 30.520 ;
        RECT 45.290 29.660 45.460 30.530 ;
        RECT 45.730 30.490 46.150 30.770 ;
        RECT 47.370 30.660 47.540 30.990 ;
        RECT 48.990 30.700 49.250 30.790 ;
        RECT 49.900 30.700 50.160 30.790 ;
        RECT 46.670 30.490 48.090 30.660 ;
        RECT 48.900 30.490 49.320 30.700 ;
        RECT 49.830 30.490 50.250 30.700 ;
        RECT 45.730 30.050 47.310 30.220 ;
        RECT 48.520 30.100 48.690 30.430 ;
        RECT 42.560 29.280 42.730 29.610 ;
        RECT 43.970 29.490 45.550 29.660 ;
        RECT 41.030 29.010 41.450 29.220 ;
        RECT 41.920 29.010 42.340 29.220 ;
        RECT 43.150 29.050 44.610 29.220 ;
        RECT 41.100 28.950 41.360 29.010 ;
        RECT 42.010 28.950 42.270 29.010 ;
        RECT 39.520 28.170 39.690 28.880 ;
        RECT 37.490 27.890 37.750 27.980 ;
        RECT 38.400 27.890 38.660 27.980 ;
        RECT 35.170 27.680 36.590 27.850 ;
        RECT 37.400 27.680 37.820 27.890 ;
        RECT 38.330 27.680 38.750 27.890 ;
        RECT 34.230 27.240 35.810 27.410 ;
        RECT 37.020 27.290 37.190 27.620 ;
        RECT 31.060 26.470 31.230 26.800 ;
        RECT 32.470 26.680 34.050 26.850 ;
        RECT 29.530 26.200 29.950 26.410 ;
        RECT 30.420 26.200 30.840 26.410 ;
        RECT 31.650 26.240 33.110 26.410 ;
        RECT 29.600 26.140 29.860 26.200 ;
        RECT 30.510 26.140 30.770 26.200 ;
        RECT 32.110 26.180 32.400 26.240 ;
        RECT 33.630 26.070 34.050 26.410 ;
        RECT 34.310 26.370 34.480 27.240 ;
        RECT 34.860 26.370 35.030 27.060 ;
        RECT 39.000 27.020 39.170 27.710 ;
        RECT 39.540 26.850 39.710 27.720 ;
        RECT 39.980 27.680 40.400 27.960 ;
        RECT 41.620 27.850 41.790 28.260 ;
        RECT 43.270 28.170 43.440 29.050 ;
        RECT 43.610 28.990 43.900 29.050 ;
        RECT 45.130 28.880 45.550 29.220 ;
        RECT 45.810 29.180 45.980 30.050 ;
        RECT 46.360 29.180 46.530 29.870 ;
        RECT 50.500 29.830 50.670 30.520 ;
        RECT 51.040 29.660 51.210 30.530 ;
        RECT 51.480 30.490 51.900 30.770 ;
        RECT 53.120 30.660 53.290 30.990 ;
        RECT 54.740 30.700 55.000 30.790 ;
        RECT 55.650 30.700 55.910 30.790 ;
        RECT 52.420 30.490 53.840 30.660 ;
        RECT 54.650 30.490 55.070 30.700 ;
        RECT 55.580 30.490 56.000 30.700 ;
        RECT 51.480 30.050 53.060 30.220 ;
        RECT 54.270 30.100 54.440 30.430 ;
        RECT 48.310 29.280 48.480 29.610 ;
        RECT 49.720 29.490 51.300 29.660 ;
        RECT 46.780 29.010 47.200 29.220 ;
        RECT 47.670 29.010 48.090 29.220 ;
        RECT 48.900 29.050 50.360 29.220 ;
        RECT 46.850 28.950 47.110 29.010 ;
        RECT 47.760 28.950 48.020 29.010 ;
        RECT 45.270 28.170 45.440 28.880 ;
        RECT 43.240 27.890 43.500 27.980 ;
        RECT 44.150 27.890 44.410 27.980 ;
        RECT 40.920 27.680 42.340 27.850 ;
        RECT 43.150 27.680 43.570 27.890 ;
        RECT 44.080 27.680 44.500 27.890 ;
        RECT 39.980 27.240 41.560 27.410 ;
        RECT 42.770 27.290 42.940 27.620 ;
        RECT 36.810 26.470 36.980 26.800 ;
        RECT 38.220 26.680 39.800 26.850 ;
        RECT 35.280 26.200 35.700 26.410 ;
        RECT 36.170 26.200 36.590 26.410 ;
        RECT 37.400 26.240 38.860 26.410 ;
        RECT 35.350 26.140 35.610 26.200 ;
        RECT 36.260 26.140 36.520 26.200 ;
        RECT 37.860 26.180 38.150 26.240 ;
        RECT 39.380 26.070 39.800 26.410 ;
        RECT 40.060 26.370 40.230 27.240 ;
        RECT 40.610 26.370 40.780 27.060 ;
        RECT 44.750 27.020 44.920 27.710 ;
        RECT 45.290 26.850 45.460 27.720 ;
        RECT 45.730 27.680 46.150 27.960 ;
        RECT 47.370 27.850 47.540 28.260 ;
        RECT 49.020 28.170 49.190 29.050 ;
        RECT 49.360 28.990 49.650 29.050 ;
        RECT 50.880 28.880 51.300 29.220 ;
        RECT 51.560 29.180 51.730 30.050 ;
        RECT 52.110 29.180 52.280 29.870 ;
        RECT 56.250 29.830 56.420 30.520 ;
        RECT 56.790 29.660 56.960 30.530 ;
        RECT 57.230 30.490 57.650 30.770 ;
        RECT 58.870 30.660 59.040 30.990 ;
        RECT 60.490 30.700 60.750 30.790 ;
        RECT 61.400 30.700 61.660 30.790 ;
        RECT 58.170 30.490 59.590 30.660 ;
        RECT 60.400 30.490 60.820 30.700 ;
        RECT 61.330 30.490 61.750 30.700 ;
        RECT 57.230 30.050 58.810 30.220 ;
        RECT 60.020 30.100 60.190 30.430 ;
        RECT 54.060 29.280 54.230 29.610 ;
        RECT 55.470 29.490 57.050 29.660 ;
        RECT 52.530 29.010 52.950 29.220 ;
        RECT 53.420 29.010 53.840 29.220 ;
        RECT 54.650 29.050 56.110 29.220 ;
        RECT 52.600 28.950 52.860 29.010 ;
        RECT 53.510 28.950 53.770 29.010 ;
        RECT 51.020 28.170 51.190 28.880 ;
        RECT 48.990 27.890 49.250 27.980 ;
        RECT 49.900 27.890 50.160 27.980 ;
        RECT 46.670 27.680 48.090 27.850 ;
        RECT 48.900 27.680 49.320 27.890 ;
        RECT 49.830 27.680 50.250 27.890 ;
        RECT 45.730 27.240 47.310 27.410 ;
        RECT 48.520 27.290 48.690 27.620 ;
        RECT 42.560 26.470 42.730 26.800 ;
        RECT 43.970 26.680 45.550 26.850 ;
        RECT 41.030 26.200 41.450 26.410 ;
        RECT 41.920 26.200 42.340 26.410 ;
        RECT 43.150 26.240 44.610 26.410 ;
        RECT 41.100 26.140 41.360 26.200 ;
        RECT 42.010 26.140 42.270 26.200 ;
        RECT 43.610 26.180 43.900 26.240 ;
        RECT 45.130 26.070 45.550 26.410 ;
        RECT 45.810 26.370 45.980 27.240 ;
        RECT 46.360 26.370 46.530 27.060 ;
        RECT 50.500 27.020 50.670 27.710 ;
        RECT 51.040 26.850 51.210 27.720 ;
        RECT 51.480 27.680 51.900 27.960 ;
        RECT 53.120 27.850 53.290 28.260 ;
        RECT 54.770 28.170 54.940 29.050 ;
        RECT 55.110 28.990 55.400 29.050 ;
        RECT 56.630 28.880 57.050 29.220 ;
        RECT 57.310 29.180 57.480 30.050 ;
        RECT 57.860 29.180 58.030 29.870 ;
        RECT 62.000 29.830 62.170 30.520 ;
        RECT 62.540 29.660 62.710 30.530 ;
        RECT 62.980 30.490 63.400 30.770 ;
        RECT 64.620 30.660 64.790 30.990 ;
        RECT 66.240 30.700 66.500 30.790 ;
        RECT 67.150 30.700 67.410 30.790 ;
        RECT 63.920 30.490 65.340 30.660 ;
        RECT 66.150 30.490 66.570 30.700 ;
        RECT 67.080 30.490 67.500 30.700 ;
        RECT 62.980 30.050 64.560 30.220 ;
        RECT 65.770 30.100 65.940 30.430 ;
        RECT 59.810 29.280 59.980 29.610 ;
        RECT 61.220 29.490 62.800 29.660 ;
        RECT 58.280 29.010 58.700 29.220 ;
        RECT 59.170 29.010 59.590 29.220 ;
        RECT 60.400 29.050 61.860 29.220 ;
        RECT 58.350 28.950 58.610 29.010 ;
        RECT 59.260 28.950 59.520 29.010 ;
        RECT 56.770 28.170 56.940 28.880 ;
        RECT 54.740 27.890 55.000 27.980 ;
        RECT 55.650 27.890 55.910 27.980 ;
        RECT 52.420 27.680 53.840 27.850 ;
        RECT 54.650 27.680 55.070 27.890 ;
        RECT 55.580 27.680 56.000 27.890 ;
        RECT 51.480 27.240 53.060 27.410 ;
        RECT 54.270 27.290 54.440 27.620 ;
        RECT 48.310 26.470 48.480 26.800 ;
        RECT 49.720 26.680 51.300 26.850 ;
        RECT 46.780 26.200 47.200 26.410 ;
        RECT 47.670 26.200 48.090 26.410 ;
        RECT 48.900 26.240 50.360 26.410 ;
        RECT 46.850 26.140 47.110 26.200 ;
        RECT 47.760 26.140 48.020 26.200 ;
        RECT 49.360 26.180 49.650 26.240 ;
        RECT 50.880 26.070 51.300 26.410 ;
        RECT 51.560 26.370 51.730 27.240 ;
        RECT 52.110 26.370 52.280 27.060 ;
        RECT 56.250 27.020 56.420 27.710 ;
        RECT 56.790 26.850 56.960 27.720 ;
        RECT 57.230 27.680 57.650 27.960 ;
        RECT 58.870 27.850 59.040 28.260 ;
        RECT 60.520 28.170 60.690 29.050 ;
        RECT 60.860 28.990 61.150 29.050 ;
        RECT 62.380 28.880 62.800 29.220 ;
        RECT 63.060 29.180 63.230 30.050 ;
        RECT 63.610 29.180 63.780 29.870 ;
        RECT 67.750 29.830 67.920 30.520 ;
        RECT 68.290 29.660 68.460 30.530 ;
        RECT 68.730 30.490 69.150 30.770 ;
        RECT 70.370 30.660 70.540 30.990 ;
        RECT 71.990 30.700 72.250 30.790 ;
        RECT 72.900 30.700 73.160 30.790 ;
        RECT 69.670 30.490 71.090 30.660 ;
        RECT 71.900 30.490 72.320 30.700 ;
        RECT 72.830 30.490 73.250 30.700 ;
        RECT 68.730 30.050 70.310 30.220 ;
        RECT 71.520 30.100 71.690 30.430 ;
        RECT 65.560 29.280 65.730 29.610 ;
        RECT 66.970 29.490 68.550 29.660 ;
        RECT 64.030 29.010 64.450 29.220 ;
        RECT 64.920 29.010 65.340 29.220 ;
        RECT 66.150 29.050 67.610 29.220 ;
        RECT 64.100 28.950 64.360 29.010 ;
        RECT 65.010 28.950 65.270 29.010 ;
        RECT 62.520 28.170 62.690 28.880 ;
        RECT 60.490 27.890 60.750 27.980 ;
        RECT 61.400 27.890 61.660 27.980 ;
        RECT 58.170 27.680 59.590 27.850 ;
        RECT 60.400 27.680 60.820 27.890 ;
        RECT 61.330 27.680 61.750 27.890 ;
        RECT 57.230 27.240 58.810 27.410 ;
        RECT 60.020 27.290 60.190 27.620 ;
        RECT 54.060 26.470 54.230 26.800 ;
        RECT 55.470 26.680 57.050 26.850 ;
        RECT 52.530 26.200 52.950 26.410 ;
        RECT 53.420 26.200 53.840 26.410 ;
        RECT 54.650 26.240 56.110 26.410 ;
        RECT 52.600 26.140 52.860 26.200 ;
        RECT 53.510 26.140 53.770 26.200 ;
        RECT 55.110 26.180 55.400 26.240 ;
        RECT 56.630 26.070 57.050 26.410 ;
        RECT 57.310 26.370 57.480 27.240 ;
        RECT 57.860 26.370 58.030 27.060 ;
        RECT 62.000 27.020 62.170 27.710 ;
        RECT 62.540 26.850 62.710 27.720 ;
        RECT 62.980 27.680 63.400 27.960 ;
        RECT 64.620 27.850 64.790 28.260 ;
        RECT 66.270 28.170 66.440 29.050 ;
        RECT 66.610 28.990 66.900 29.050 ;
        RECT 68.130 28.880 68.550 29.220 ;
        RECT 68.810 29.180 68.980 30.050 ;
        RECT 69.360 29.180 69.530 29.870 ;
        RECT 73.500 29.830 73.670 30.520 ;
        RECT 74.040 29.660 74.210 30.530 ;
        RECT 74.480 30.490 74.900 30.770 ;
        RECT 76.120 30.660 76.290 30.990 ;
        RECT 77.740 30.700 78.000 30.790 ;
        RECT 78.650 30.700 78.910 30.790 ;
        RECT 75.420 30.490 76.840 30.660 ;
        RECT 77.650 30.490 78.070 30.700 ;
        RECT 78.580 30.490 79.000 30.700 ;
        RECT 74.480 30.050 76.060 30.220 ;
        RECT 77.270 30.100 77.440 30.430 ;
        RECT 71.310 29.280 71.480 29.610 ;
        RECT 72.720 29.490 74.300 29.660 ;
        RECT 69.780 29.010 70.200 29.220 ;
        RECT 70.670 29.010 71.090 29.220 ;
        RECT 71.900 29.050 73.360 29.220 ;
        RECT 69.850 28.950 70.110 29.010 ;
        RECT 70.760 28.950 71.020 29.010 ;
        RECT 68.270 28.170 68.440 28.880 ;
        RECT 66.240 27.890 66.500 27.980 ;
        RECT 67.150 27.890 67.410 27.980 ;
        RECT 63.920 27.680 65.340 27.850 ;
        RECT 66.150 27.680 66.570 27.890 ;
        RECT 67.080 27.680 67.500 27.890 ;
        RECT 62.980 27.240 64.560 27.410 ;
        RECT 65.770 27.290 65.940 27.620 ;
        RECT 59.810 26.470 59.980 26.800 ;
        RECT 61.220 26.680 62.800 26.850 ;
        RECT 58.280 26.200 58.700 26.410 ;
        RECT 59.170 26.200 59.590 26.410 ;
        RECT 60.400 26.240 61.860 26.410 ;
        RECT 58.350 26.140 58.610 26.200 ;
        RECT 59.260 26.140 59.520 26.200 ;
        RECT 60.860 26.180 61.150 26.240 ;
        RECT 62.380 26.070 62.800 26.410 ;
        RECT 63.060 26.370 63.230 27.240 ;
        RECT 63.610 26.370 63.780 27.060 ;
        RECT 67.750 27.020 67.920 27.710 ;
        RECT 68.290 26.850 68.460 27.720 ;
        RECT 68.730 27.680 69.150 27.960 ;
        RECT 70.370 27.850 70.540 28.260 ;
        RECT 72.020 28.170 72.190 29.050 ;
        RECT 72.360 28.990 72.650 29.050 ;
        RECT 73.880 28.880 74.300 29.220 ;
        RECT 74.560 29.180 74.730 30.050 ;
        RECT 75.110 29.180 75.280 29.870 ;
        RECT 79.250 29.830 79.420 30.520 ;
        RECT 79.790 29.660 79.960 30.530 ;
        RECT 80.230 30.490 80.650 30.770 ;
        RECT 81.870 30.660 82.040 30.990 ;
        RECT 83.490 30.700 83.750 30.790 ;
        RECT 84.400 30.700 84.660 30.790 ;
        RECT 81.170 30.490 82.590 30.660 ;
        RECT 83.400 30.490 83.820 30.700 ;
        RECT 84.330 30.490 84.750 30.700 ;
        RECT 80.230 30.050 81.810 30.220 ;
        RECT 83.020 30.100 83.190 30.430 ;
        RECT 77.060 29.280 77.230 29.610 ;
        RECT 78.470 29.490 80.050 29.660 ;
        RECT 75.530 29.010 75.950 29.220 ;
        RECT 76.420 29.010 76.840 29.220 ;
        RECT 77.650 29.050 79.110 29.220 ;
        RECT 75.600 28.950 75.860 29.010 ;
        RECT 76.510 28.950 76.770 29.010 ;
        RECT 74.020 28.170 74.190 28.880 ;
        RECT 71.990 27.890 72.250 27.980 ;
        RECT 72.900 27.890 73.160 27.980 ;
        RECT 69.670 27.680 71.090 27.850 ;
        RECT 71.900 27.680 72.320 27.890 ;
        RECT 72.830 27.680 73.250 27.890 ;
        RECT 68.730 27.240 70.310 27.410 ;
        RECT 71.520 27.290 71.690 27.620 ;
        RECT 65.560 26.470 65.730 26.800 ;
        RECT 66.970 26.680 68.550 26.850 ;
        RECT 64.030 26.200 64.450 26.410 ;
        RECT 64.920 26.200 65.340 26.410 ;
        RECT 66.150 26.240 67.610 26.410 ;
        RECT 64.100 26.140 64.360 26.200 ;
        RECT 65.010 26.140 65.270 26.200 ;
        RECT 66.610 26.180 66.900 26.240 ;
        RECT 68.130 26.070 68.550 26.410 ;
        RECT 68.810 26.370 68.980 27.240 ;
        RECT 69.360 26.370 69.530 27.060 ;
        RECT 73.500 27.020 73.670 27.710 ;
        RECT 74.040 26.850 74.210 27.720 ;
        RECT 74.480 27.680 74.900 27.960 ;
        RECT 76.120 27.850 76.290 28.260 ;
        RECT 77.770 28.170 77.940 29.050 ;
        RECT 78.110 28.990 78.400 29.050 ;
        RECT 79.630 28.880 80.050 29.220 ;
        RECT 80.310 29.180 80.480 30.050 ;
        RECT 80.860 29.180 81.030 29.870 ;
        RECT 85.000 29.830 85.170 30.520 ;
        RECT 85.540 29.660 85.710 30.530 ;
        RECT 85.980 30.490 86.400 30.770 ;
        RECT 87.620 30.660 87.790 30.990 ;
        RECT 89.240 30.700 89.500 30.790 ;
        RECT 90.150 30.700 90.410 30.790 ;
        RECT 86.920 30.490 88.340 30.660 ;
        RECT 89.150 30.490 89.570 30.700 ;
        RECT 90.080 30.490 90.500 30.700 ;
        RECT 85.980 30.050 87.560 30.220 ;
        RECT 88.770 30.100 88.940 30.430 ;
        RECT 82.810 29.280 82.980 29.610 ;
        RECT 84.220 29.490 85.800 29.660 ;
        RECT 81.280 29.010 81.700 29.220 ;
        RECT 82.170 29.010 82.590 29.220 ;
        RECT 83.400 29.050 84.860 29.220 ;
        RECT 81.350 28.950 81.610 29.010 ;
        RECT 82.260 28.950 82.520 29.010 ;
        RECT 79.770 28.170 79.940 28.880 ;
        RECT 77.740 27.890 78.000 27.980 ;
        RECT 78.650 27.890 78.910 27.980 ;
        RECT 75.420 27.680 76.840 27.850 ;
        RECT 77.650 27.680 78.070 27.890 ;
        RECT 78.580 27.680 79.000 27.890 ;
        RECT 74.480 27.240 76.060 27.410 ;
        RECT 77.270 27.290 77.440 27.620 ;
        RECT 71.310 26.470 71.480 26.800 ;
        RECT 72.720 26.680 74.300 26.850 ;
        RECT 69.780 26.200 70.200 26.410 ;
        RECT 70.670 26.200 71.090 26.410 ;
        RECT 71.900 26.240 73.360 26.410 ;
        RECT 69.850 26.140 70.110 26.200 ;
        RECT 70.760 26.140 71.020 26.200 ;
        RECT 72.360 26.180 72.650 26.240 ;
        RECT 73.880 26.070 74.300 26.410 ;
        RECT 74.560 26.370 74.730 27.240 ;
        RECT 75.110 26.370 75.280 27.060 ;
        RECT 79.250 27.020 79.420 27.710 ;
        RECT 79.790 26.850 79.960 27.720 ;
        RECT 80.230 27.680 80.650 27.960 ;
        RECT 81.870 27.850 82.040 28.260 ;
        RECT 83.520 28.170 83.690 29.050 ;
        RECT 83.860 28.990 84.150 29.050 ;
        RECT 85.380 28.880 85.800 29.220 ;
        RECT 86.060 29.180 86.230 30.050 ;
        RECT 86.610 29.180 86.780 29.870 ;
        RECT 90.750 29.830 90.920 30.520 ;
        RECT 91.290 29.660 91.460 30.530 ;
        RECT 91.730 30.490 92.150 30.770 ;
        RECT 93.370 30.660 93.540 30.990 ;
        RECT 92.670 30.490 94.090 30.660 ;
        RECT 91.730 30.050 93.310 30.220 ;
        RECT 88.560 29.280 88.730 29.610 ;
        RECT 89.970 29.490 91.550 29.660 ;
        RECT 87.030 29.010 87.450 29.220 ;
        RECT 87.920 29.010 88.340 29.220 ;
        RECT 89.150 29.050 90.610 29.220 ;
        RECT 87.100 28.950 87.360 29.010 ;
        RECT 88.010 28.950 88.270 29.010 ;
        RECT 85.520 28.170 85.690 28.880 ;
        RECT 83.490 27.890 83.750 27.980 ;
        RECT 84.400 27.890 84.660 27.980 ;
        RECT 81.170 27.680 82.590 27.850 ;
        RECT 83.400 27.680 83.820 27.890 ;
        RECT 84.330 27.680 84.750 27.890 ;
        RECT 80.230 27.240 81.810 27.410 ;
        RECT 83.020 27.290 83.190 27.620 ;
        RECT 77.060 26.470 77.230 26.800 ;
        RECT 78.470 26.680 80.050 26.850 ;
        RECT 75.530 26.200 75.950 26.410 ;
        RECT 76.420 26.200 76.840 26.410 ;
        RECT 77.650 26.240 79.110 26.410 ;
        RECT 75.600 26.140 75.860 26.200 ;
        RECT 76.510 26.140 76.770 26.200 ;
        RECT 78.110 26.180 78.400 26.240 ;
        RECT 79.630 26.070 80.050 26.410 ;
        RECT 80.310 26.370 80.480 27.240 ;
        RECT 80.860 26.370 81.030 27.060 ;
        RECT 85.000 27.020 85.170 27.710 ;
        RECT 85.540 26.850 85.710 27.720 ;
        RECT 85.980 27.680 86.400 27.960 ;
        RECT 87.620 27.850 87.790 28.260 ;
        RECT 89.270 28.170 89.440 29.050 ;
        RECT 89.610 28.990 89.900 29.050 ;
        RECT 91.130 28.880 91.550 29.220 ;
        RECT 91.810 29.180 91.980 30.050 ;
        RECT 92.360 29.180 92.530 29.870 ;
        RECT 94.310 29.280 94.480 29.610 ;
        RECT 92.780 29.010 93.200 29.220 ;
        RECT 93.670 29.010 94.090 29.220 ;
        RECT 92.850 28.950 93.110 29.010 ;
        RECT 93.760 28.950 94.020 29.010 ;
        RECT 91.270 28.170 91.440 28.880 ;
        RECT 94.230 28.260 94.400 28.530 ;
        RECT 93.370 28.090 94.400 28.260 ;
        RECT 89.240 27.890 89.500 27.980 ;
        RECT 90.150 27.890 90.410 27.980 ;
        RECT 86.920 27.680 88.340 27.850 ;
        RECT 89.150 27.680 89.570 27.890 ;
        RECT 90.080 27.680 90.500 27.890 ;
        RECT 85.980 27.240 87.560 27.410 ;
        RECT 88.770 27.290 88.940 27.620 ;
        RECT 82.810 26.470 82.980 26.800 ;
        RECT 84.220 26.680 85.800 26.850 ;
        RECT 81.280 26.200 81.700 26.410 ;
        RECT 82.170 26.200 82.590 26.410 ;
        RECT 83.400 26.240 84.860 26.410 ;
        RECT 81.350 26.140 81.610 26.200 ;
        RECT 82.260 26.140 82.520 26.200 ;
        RECT 83.860 26.180 84.150 26.240 ;
        RECT 85.380 26.070 85.800 26.410 ;
        RECT 86.060 26.370 86.230 27.240 ;
        RECT 86.610 26.370 86.780 27.060 ;
        RECT 90.750 27.020 90.920 27.710 ;
        RECT 91.290 26.850 91.460 27.720 ;
        RECT 91.730 27.680 92.150 27.960 ;
        RECT 93.370 27.850 93.540 28.090 ;
        RECT 92.670 27.680 94.090 27.850 ;
        RECT 91.730 27.240 93.310 27.410 ;
        RECT 88.560 26.470 88.730 26.800 ;
        RECT 89.970 26.680 91.550 26.850 ;
        RECT 87.030 26.200 87.450 26.410 ;
        RECT 87.920 26.200 88.340 26.410 ;
        RECT 89.150 26.240 90.610 26.410 ;
        RECT 87.100 26.140 87.360 26.200 ;
        RECT 88.010 26.140 88.270 26.200 ;
        RECT 89.610 26.180 89.900 26.240 ;
        RECT 91.130 26.070 91.550 26.410 ;
        RECT 91.810 26.370 91.980 27.240 ;
        RECT 92.360 26.370 92.530 27.060 ;
        RECT 94.310 26.470 94.480 26.800 ;
        RECT 92.780 26.200 93.200 26.410 ;
        RECT 93.670 26.200 94.090 26.410 ;
        RECT 92.850 26.140 93.110 26.200 ;
        RECT 93.760 26.140 94.020 26.200 ;
        RECT 2.990 25.480 3.250 25.570 ;
        RECT 3.900 25.480 4.160 25.570 ;
        RECT 2.900 25.270 3.320 25.480 ;
        RECT 3.830 25.270 4.250 25.480 ;
        RECT 2.520 24.880 2.690 25.210 ;
        RECT 4.500 24.610 4.670 25.300 ;
        RECT 5.040 24.440 5.210 25.310 ;
        RECT 5.480 25.270 5.900 25.550 ;
        RECT 7.120 25.440 7.290 25.770 ;
        RECT 8.740 25.480 9.000 25.570 ;
        RECT 9.650 25.480 9.910 25.570 ;
        RECT 6.420 25.270 7.840 25.440 ;
        RECT 8.650 25.270 9.070 25.480 ;
        RECT 9.580 25.270 10.000 25.480 ;
        RECT 5.480 24.830 7.060 25.000 ;
        RECT 8.270 24.880 8.440 25.210 ;
        RECT 3.720 24.270 5.300 24.440 ;
        RECT 2.900 23.830 4.360 24.000 ;
        RECT 3.360 23.770 3.650 23.830 ;
        RECT 4.880 23.660 5.300 24.000 ;
        RECT 5.560 23.960 5.730 24.830 ;
        RECT 6.110 23.960 6.280 24.650 ;
        RECT 10.250 24.610 10.420 25.300 ;
        RECT 10.790 24.440 10.960 25.310 ;
        RECT 11.230 25.270 11.650 25.550 ;
        RECT 12.870 25.440 13.040 25.770 ;
        RECT 14.490 25.480 14.750 25.570 ;
        RECT 15.400 25.480 15.660 25.570 ;
        RECT 12.170 25.270 13.590 25.440 ;
        RECT 14.400 25.270 14.820 25.480 ;
        RECT 15.330 25.270 15.750 25.480 ;
        RECT 11.230 24.830 12.810 25.000 ;
        RECT 14.020 24.880 14.190 25.210 ;
        RECT 8.060 24.060 8.230 24.390 ;
        RECT 9.470 24.270 11.050 24.440 ;
        RECT 6.530 23.790 6.950 24.000 ;
        RECT 7.420 23.790 7.840 24.000 ;
        RECT 8.650 23.830 10.110 24.000 ;
        RECT 6.600 23.730 6.860 23.790 ;
        RECT 7.510 23.730 7.770 23.790 ;
        RECT 9.110 23.770 9.400 23.830 ;
        RECT 10.630 23.660 11.050 24.000 ;
        RECT 11.310 23.960 11.480 24.830 ;
        RECT 11.860 23.960 12.030 24.650 ;
        RECT 16.000 24.610 16.170 25.300 ;
        RECT 16.540 24.440 16.710 25.310 ;
        RECT 16.980 25.270 17.400 25.550 ;
        RECT 18.620 25.440 18.790 25.770 ;
        RECT 20.240 25.480 20.500 25.570 ;
        RECT 21.150 25.480 21.410 25.570 ;
        RECT 17.920 25.270 19.340 25.440 ;
        RECT 20.150 25.270 20.570 25.480 ;
        RECT 21.080 25.270 21.500 25.480 ;
        RECT 16.980 24.830 18.560 25.000 ;
        RECT 19.770 24.880 19.940 25.210 ;
        RECT 13.810 24.060 13.980 24.390 ;
        RECT 15.220 24.270 16.800 24.440 ;
        RECT 12.280 23.790 12.700 24.000 ;
        RECT 13.170 23.790 13.590 24.000 ;
        RECT 14.400 23.830 15.860 24.000 ;
        RECT 12.350 23.730 12.610 23.790 ;
        RECT 13.260 23.730 13.520 23.790 ;
        RECT 14.860 23.770 15.150 23.830 ;
        RECT 16.380 23.660 16.800 24.000 ;
        RECT 17.060 23.960 17.230 24.830 ;
        RECT 17.610 23.960 17.780 24.650 ;
        RECT 21.750 24.610 21.920 25.300 ;
        RECT 22.290 24.440 22.460 25.310 ;
        RECT 22.730 25.270 23.150 25.550 ;
        RECT 24.370 25.440 24.540 25.770 ;
        RECT 25.990 25.480 26.250 25.570 ;
        RECT 26.900 25.480 27.160 25.570 ;
        RECT 23.670 25.270 25.090 25.440 ;
        RECT 25.900 25.270 26.320 25.480 ;
        RECT 26.830 25.270 27.250 25.480 ;
        RECT 22.730 24.830 24.310 25.000 ;
        RECT 25.520 24.880 25.690 25.210 ;
        RECT 19.560 24.060 19.730 24.390 ;
        RECT 20.970 24.270 22.550 24.440 ;
        RECT 18.030 23.790 18.450 24.000 ;
        RECT 18.920 23.790 19.340 24.000 ;
        RECT 20.150 23.830 21.610 24.000 ;
        RECT 18.100 23.730 18.360 23.790 ;
        RECT 19.010 23.730 19.270 23.790 ;
        RECT 20.610 23.770 20.900 23.830 ;
        RECT 22.130 23.660 22.550 24.000 ;
        RECT 22.810 23.960 22.980 24.830 ;
        RECT 23.360 23.960 23.530 24.650 ;
        RECT 27.500 24.610 27.670 25.300 ;
        RECT 28.040 24.440 28.210 25.310 ;
        RECT 28.480 25.270 28.900 25.550 ;
        RECT 30.120 25.440 30.290 25.770 ;
        RECT 31.740 25.480 32.000 25.570 ;
        RECT 32.650 25.480 32.910 25.570 ;
        RECT 29.420 25.270 30.840 25.440 ;
        RECT 31.650 25.270 32.070 25.480 ;
        RECT 32.580 25.270 33.000 25.480 ;
        RECT 28.480 24.830 30.060 25.000 ;
        RECT 31.270 24.880 31.440 25.210 ;
        RECT 25.310 24.060 25.480 24.390 ;
        RECT 26.720 24.270 28.300 24.440 ;
        RECT 23.780 23.790 24.200 24.000 ;
        RECT 24.670 23.790 25.090 24.000 ;
        RECT 25.900 23.830 27.360 24.000 ;
        RECT 23.850 23.730 24.110 23.790 ;
        RECT 24.760 23.730 25.020 23.790 ;
        RECT 26.360 23.770 26.650 23.830 ;
        RECT 27.880 23.660 28.300 24.000 ;
        RECT 28.560 23.960 28.730 24.830 ;
        RECT 29.110 23.960 29.280 24.650 ;
        RECT 33.250 24.610 33.420 25.300 ;
        RECT 33.790 24.440 33.960 25.310 ;
        RECT 34.230 25.270 34.650 25.550 ;
        RECT 35.870 25.440 36.040 25.770 ;
        RECT 37.490 25.480 37.750 25.570 ;
        RECT 38.400 25.480 38.660 25.570 ;
        RECT 35.170 25.270 36.590 25.440 ;
        RECT 37.400 25.270 37.820 25.480 ;
        RECT 38.330 25.270 38.750 25.480 ;
        RECT 34.230 24.830 35.810 25.000 ;
        RECT 37.020 24.880 37.190 25.210 ;
        RECT 31.060 24.060 31.230 24.390 ;
        RECT 32.470 24.270 34.050 24.440 ;
        RECT 29.530 23.790 29.950 24.000 ;
        RECT 30.420 23.790 30.840 24.000 ;
        RECT 31.650 23.830 33.110 24.000 ;
        RECT 29.600 23.730 29.860 23.790 ;
        RECT 30.510 23.730 30.770 23.790 ;
        RECT 32.110 23.770 32.400 23.830 ;
        RECT 33.630 23.660 34.050 24.000 ;
        RECT 34.310 23.960 34.480 24.830 ;
        RECT 34.860 23.960 35.030 24.650 ;
        RECT 39.000 24.610 39.170 25.300 ;
        RECT 39.540 24.440 39.710 25.310 ;
        RECT 39.980 25.270 40.400 25.550 ;
        RECT 41.620 25.440 41.790 25.770 ;
        RECT 43.240 25.480 43.500 25.570 ;
        RECT 44.150 25.480 44.410 25.570 ;
        RECT 40.920 25.270 42.340 25.440 ;
        RECT 43.150 25.270 43.570 25.480 ;
        RECT 44.080 25.270 44.500 25.480 ;
        RECT 39.980 24.830 41.560 25.000 ;
        RECT 42.770 24.880 42.940 25.210 ;
        RECT 36.810 24.060 36.980 24.390 ;
        RECT 38.220 24.270 39.800 24.440 ;
        RECT 35.280 23.790 35.700 24.000 ;
        RECT 36.170 23.790 36.590 24.000 ;
        RECT 37.400 23.830 38.860 24.000 ;
        RECT 35.350 23.730 35.610 23.790 ;
        RECT 36.260 23.730 36.520 23.790 ;
        RECT 37.860 23.770 38.150 23.830 ;
        RECT 39.380 23.660 39.800 24.000 ;
        RECT 40.060 23.960 40.230 24.830 ;
        RECT 40.610 23.960 40.780 24.650 ;
        RECT 44.750 24.610 44.920 25.300 ;
        RECT 45.290 24.440 45.460 25.310 ;
        RECT 45.730 25.270 46.150 25.550 ;
        RECT 47.370 25.440 47.540 25.770 ;
        RECT 48.990 25.480 49.250 25.570 ;
        RECT 49.900 25.480 50.160 25.570 ;
        RECT 46.670 25.270 48.090 25.440 ;
        RECT 48.900 25.270 49.320 25.480 ;
        RECT 49.830 25.270 50.250 25.480 ;
        RECT 45.730 24.830 47.310 25.000 ;
        RECT 48.520 24.880 48.690 25.210 ;
        RECT 42.560 24.060 42.730 24.390 ;
        RECT 43.970 24.270 45.550 24.440 ;
        RECT 41.030 23.790 41.450 24.000 ;
        RECT 41.920 23.790 42.340 24.000 ;
        RECT 43.150 23.830 44.610 24.000 ;
        RECT 41.100 23.730 41.360 23.790 ;
        RECT 42.010 23.730 42.270 23.790 ;
        RECT 43.610 23.770 43.900 23.830 ;
        RECT 45.130 23.660 45.550 24.000 ;
        RECT 45.810 23.960 45.980 24.830 ;
        RECT 46.360 23.960 46.530 24.650 ;
        RECT 50.500 24.610 50.670 25.300 ;
        RECT 51.040 24.440 51.210 25.310 ;
        RECT 51.480 25.270 51.900 25.550 ;
        RECT 53.120 25.440 53.290 25.770 ;
        RECT 54.740 25.480 55.000 25.570 ;
        RECT 55.650 25.480 55.910 25.570 ;
        RECT 52.420 25.270 53.840 25.440 ;
        RECT 54.650 25.270 55.070 25.480 ;
        RECT 55.580 25.270 56.000 25.480 ;
        RECT 51.480 24.830 53.060 25.000 ;
        RECT 54.270 24.880 54.440 25.210 ;
        RECT 48.310 24.060 48.480 24.390 ;
        RECT 49.720 24.270 51.300 24.440 ;
        RECT 46.780 23.790 47.200 24.000 ;
        RECT 47.670 23.790 48.090 24.000 ;
        RECT 48.900 23.830 50.360 24.000 ;
        RECT 46.850 23.730 47.110 23.790 ;
        RECT 47.760 23.730 48.020 23.790 ;
        RECT 49.360 23.770 49.650 23.830 ;
        RECT 50.880 23.660 51.300 24.000 ;
        RECT 51.560 23.960 51.730 24.830 ;
        RECT 52.110 23.960 52.280 24.650 ;
        RECT 56.250 24.610 56.420 25.300 ;
        RECT 56.790 24.440 56.960 25.310 ;
        RECT 57.230 25.270 57.650 25.550 ;
        RECT 58.870 25.440 59.040 25.770 ;
        RECT 60.490 25.480 60.750 25.570 ;
        RECT 61.400 25.480 61.660 25.570 ;
        RECT 58.170 25.270 59.590 25.440 ;
        RECT 60.400 25.270 60.820 25.480 ;
        RECT 61.330 25.270 61.750 25.480 ;
        RECT 57.230 24.830 58.810 25.000 ;
        RECT 60.020 24.880 60.190 25.210 ;
        RECT 54.060 24.060 54.230 24.390 ;
        RECT 55.470 24.270 57.050 24.440 ;
        RECT 52.530 23.790 52.950 24.000 ;
        RECT 53.420 23.790 53.840 24.000 ;
        RECT 54.650 23.830 56.110 24.000 ;
        RECT 52.600 23.730 52.860 23.790 ;
        RECT 53.510 23.730 53.770 23.790 ;
        RECT 55.110 23.770 55.400 23.830 ;
        RECT 56.630 23.660 57.050 24.000 ;
        RECT 57.310 23.960 57.480 24.830 ;
        RECT 57.860 23.960 58.030 24.650 ;
        RECT 62.000 24.610 62.170 25.300 ;
        RECT 62.540 24.440 62.710 25.310 ;
        RECT 62.980 25.270 63.400 25.550 ;
        RECT 64.620 25.440 64.790 25.770 ;
        RECT 66.240 25.480 66.500 25.570 ;
        RECT 67.150 25.480 67.410 25.570 ;
        RECT 63.920 25.270 65.340 25.440 ;
        RECT 66.150 25.270 66.570 25.480 ;
        RECT 67.080 25.270 67.500 25.480 ;
        RECT 62.980 24.830 64.560 25.000 ;
        RECT 65.770 24.880 65.940 25.210 ;
        RECT 59.810 24.060 59.980 24.390 ;
        RECT 61.220 24.270 62.800 24.440 ;
        RECT 58.280 23.790 58.700 24.000 ;
        RECT 59.170 23.790 59.590 24.000 ;
        RECT 60.400 23.830 61.860 24.000 ;
        RECT 58.350 23.730 58.610 23.790 ;
        RECT 59.260 23.730 59.520 23.790 ;
        RECT 60.860 23.770 61.150 23.830 ;
        RECT 62.380 23.660 62.800 24.000 ;
        RECT 63.060 23.960 63.230 24.830 ;
        RECT 63.610 23.960 63.780 24.650 ;
        RECT 67.750 24.610 67.920 25.300 ;
        RECT 68.290 24.440 68.460 25.310 ;
        RECT 68.730 25.270 69.150 25.550 ;
        RECT 70.370 25.440 70.540 25.770 ;
        RECT 71.990 25.480 72.250 25.570 ;
        RECT 72.900 25.480 73.160 25.570 ;
        RECT 69.670 25.270 71.090 25.440 ;
        RECT 71.900 25.270 72.320 25.480 ;
        RECT 72.830 25.270 73.250 25.480 ;
        RECT 68.730 24.830 70.310 25.000 ;
        RECT 71.520 24.880 71.690 25.210 ;
        RECT 65.560 24.060 65.730 24.390 ;
        RECT 66.970 24.270 68.550 24.440 ;
        RECT 64.030 23.790 64.450 24.000 ;
        RECT 64.920 23.790 65.340 24.000 ;
        RECT 66.150 23.830 67.610 24.000 ;
        RECT 64.100 23.730 64.360 23.790 ;
        RECT 65.010 23.730 65.270 23.790 ;
        RECT 66.610 23.770 66.900 23.830 ;
        RECT 68.130 23.660 68.550 24.000 ;
        RECT 68.810 23.960 68.980 24.830 ;
        RECT 69.360 23.960 69.530 24.650 ;
        RECT 73.500 24.610 73.670 25.300 ;
        RECT 74.040 24.440 74.210 25.310 ;
        RECT 74.480 25.270 74.900 25.550 ;
        RECT 76.120 25.440 76.290 25.770 ;
        RECT 77.740 25.480 78.000 25.570 ;
        RECT 78.650 25.480 78.910 25.570 ;
        RECT 75.420 25.270 76.840 25.440 ;
        RECT 77.650 25.270 78.070 25.480 ;
        RECT 78.580 25.270 79.000 25.480 ;
        RECT 74.480 24.830 76.060 25.000 ;
        RECT 77.270 24.880 77.440 25.210 ;
        RECT 71.310 24.060 71.480 24.390 ;
        RECT 72.720 24.270 74.300 24.440 ;
        RECT 69.780 23.790 70.200 24.000 ;
        RECT 70.670 23.790 71.090 24.000 ;
        RECT 71.900 23.830 73.360 24.000 ;
        RECT 69.850 23.730 70.110 23.790 ;
        RECT 70.760 23.730 71.020 23.790 ;
        RECT 72.360 23.770 72.650 23.830 ;
        RECT 73.880 23.660 74.300 24.000 ;
        RECT 74.560 23.960 74.730 24.830 ;
        RECT 75.110 23.960 75.280 24.650 ;
        RECT 79.250 24.610 79.420 25.300 ;
        RECT 79.790 24.440 79.960 25.310 ;
        RECT 80.230 25.270 80.650 25.550 ;
        RECT 81.870 25.440 82.040 25.770 ;
        RECT 83.490 25.480 83.750 25.570 ;
        RECT 84.400 25.480 84.660 25.570 ;
        RECT 81.170 25.270 82.590 25.440 ;
        RECT 83.400 25.270 83.820 25.480 ;
        RECT 84.330 25.270 84.750 25.480 ;
        RECT 80.230 24.830 81.810 25.000 ;
        RECT 83.020 24.880 83.190 25.210 ;
        RECT 77.060 24.060 77.230 24.390 ;
        RECT 78.470 24.270 80.050 24.440 ;
        RECT 75.530 23.790 75.950 24.000 ;
        RECT 76.420 23.790 76.840 24.000 ;
        RECT 77.650 23.830 79.110 24.000 ;
        RECT 75.600 23.730 75.860 23.790 ;
        RECT 76.510 23.730 76.770 23.790 ;
        RECT 78.110 23.770 78.400 23.830 ;
        RECT 79.630 23.660 80.050 24.000 ;
        RECT 80.310 23.960 80.480 24.830 ;
        RECT 80.860 23.960 81.030 24.650 ;
        RECT 85.000 24.610 85.170 25.300 ;
        RECT 85.540 24.440 85.710 25.310 ;
        RECT 85.980 25.270 86.400 25.550 ;
        RECT 87.620 25.440 87.790 25.770 ;
        RECT 89.240 25.480 89.500 25.570 ;
        RECT 90.150 25.480 90.410 25.570 ;
        RECT 86.920 25.270 88.340 25.440 ;
        RECT 89.150 25.270 89.570 25.480 ;
        RECT 90.080 25.270 90.500 25.480 ;
        RECT 85.980 24.830 87.560 25.000 ;
        RECT 88.770 24.880 88.940 25.210 ;
        RECT 82.810 24.060 82.980 24.390 ;
        RECT 84.220 24.270 85.800 24.440 ;
        RECT 81.280 23.790 81.700 24.000 ;
        RECT 82.170 23.790 82.590 24.000 ;
        RECT 83.400 23.830 84.860 24.000 ;
        RECT 81.350 23.730 81.610 23.790 ;
        RECT 82.260 23.730 82.520 23.790 ;
        RECT 83.860 23.770 84.150 23.830 ;
        RECT 85.380 23.660 85.800 24.000 ;
        RECT 86.060 23.960 86.230 24.830 ;
        RECT 86.610 23.960 86.780 24.650 ;
        RECT 90.750 24.610 90.920 25.300 ;
        RECT 91.290 24.440 91.460 25.310 ;
        RECT 91.730 25.270 92.150 25.550 ;
        RECT 93.370 25.440 93.540 25.770 ;
        RECT 92.670 25.270 94.090 25.440 ;
        RECT 91.730 24.830 93.310 25.000 ;
        RECT 88.560 24.060 88.730 24.390 ;
        RECT 89.970 24.270 91.550 24.440 ;
        RECT 87.030 23.790 87.450 24.000 ;
        RECT 87.920 23.790 88.340 24.000 ;
        RECT 89.150 23.830 90.610 24.000 ;
        RECT 87.100 23.730 87.360 23.790 ;
        RECT 88.010 23.730 88.270 23.790 ;
        RECT 89.610 23.770 89.900 23.830 ;
        RECT 91.130 23.660 91.550 24.000 ;
        RECT 91.810 23.960 91.980 24.830 ;
        RECT 92.360 23.960 92.530 24.650 ;
        RECT 94.310 24.060 94.480 24.390 ;
        RECT 92.780 23.790 93.200 24.000 ;
        RECT 93.670 23.790 94.090 24.000 ;
        RECT 92.850 23.730 93.110 23.790 ;
        RECT 93.760 23.730 94.020 23.790 ;
        RECT 2.990 23.070 3.250 23.160 ;
        RECT 3.900 23.070 4.160 23.160 ;
        RECT 2.900 22.860 3.320 23.070 ;
        RECT 3.830 22.860 4.250 23.070 ;
        RECT 2.520 22.470 2.690 22.800 ;
        RECT 4.500 22.200 4.670 22.890 ;
        RECT 5.040 22.030 5.210 22.900 ;
        RECT 5.480 22.860 5.900 23.140 ;
        RECT 7.120 23.030 7.290 23.360 ;
        RECT 8.740 23.070 9.000 23.160 ;
        RECT 9.650 23.070 9.910 23.160 ;
        RECT 6.420 22.860 7.840 23.030 ;
        RECT 8.650 22.860 9.070 23.070 ;
        RECT 9.580 22.860 10.000 23.070 ;
        RECT 5.480 22.420 7.060 22.590 ;
        RECT 8.270 22.470 8.440 22.800 ;
        RECT 3.720 21.860 5.300 22.030 ;
        RECT 2.900 21.420 4.360 21.590 ;
        RECT 3.360 21.360 3.650 21.420 ;
        RECT 4.880 21.250 5.300 21.590 ;
        RECT 5.560 21.550 5.730 22.420 ;
        RECT 6.110 21.550 6.280 22.240 ;
        RECT 10.250 22.200 10.420 22.890 ;
        RECT 10.790 22.030 10.960 22.900 ;
        RECT 11.230 22.860 11.650 23.140 ;
        RECT 12.870 23.030 13.040 23.360 ;
        RECT 14.490 23.070 14.750 23.160 ;
        RECT 15.400 23.070 15.660 23.160 ;
        RECT 12.170 22.860 13.590 23.030 ;
        RECT 14.400 22.860 14.820 23.070 ;
        RECT 15.330 22.860 15.750 23.070 ;
        RECT 11.230 22.420 12.810 22.590 ;
        RECT 14.020 22.470 14.190 22.800 ;
        RECT 8.060 21.650 8.230 21.980 ;
        RECT 9.470 21.860 11.050 22.030 ;
        RECT 6.530 21.380 6.950 21.590 ;
        RECT 7.420 21.380 7.840 21.590 ;
        RECT 8.650 21.420 10.110 21.590 ;
        RECT 6.600 21.320 6.860 21.380 ;
        RECT 7.510 21.320 7.770 21.380 ;
        RECT 9.110 21.360 9.400 21.420 ;
        RECT 10.630 21.250 11.050 21.590 ;
        RECT 11.310 21.550 11.480 22.420 ;
        RECT 11.860 21.550 12.030 22.240 ;
        RECT 16.000 22.200 16.170 22.890 ;
        RECT 16.540 22.030 16.710 22.900 ;
        RECT 16.980 22.860 17.400 23.140 ;
        RECT 18.620 23.030 18.790 23.360 ;
        RECT 20.240 23.070 20.500 23.160 ;
        RECT 21.150 23.070 21.410 23.160 ;
        RECT 17.920 22.860 19.340 23.030 ;
        RECT 20.150 22.860 20.570 23.070 ;
        RECT 21.080 22.860 21.500 23.070 ;
        RECT 16.980 22.420 18.560 22.590 ;
        RECT 19.770 22.470 19.940 22.800 ;
        RECT 13.810 21.650 13.980 21.980 ;
        RECT 15.220 21.860 16.800 22.030 ;
        RECT 12.280 21.380 12.700 21.590 ;
        RECT 13.170 21.380 13.590 21.590 ;
        RECT 14.400 21.420 15.860 21.590 ;
        RECT 12.350 21.320 12.610 21.380 ;
        RECT 13.260 21.320 13.520 21.380 ;
        RECT 14.860 21.360 15.150 21.420 ;
        RECT 16.380 21.250 16.800 21.590 ;
        RECT 17.060 21.550 17.230 22.420 ;
        RECT 17.610 21.550 17.780 22.240 ;
        RECT 21.750 22.200 21.920 22.890 ;
        RECT 22.290 22.030 22.460 22.900 ;
        RECT 22.730 22.860 23.150 23.140 ;
        RECT 24.370 23.030 24.540 23.360 ;
        RECT 25.990 23.070 26.250 23.160 ;
        RECT 26.900 23.070 27.160 23.160 ;
        RECT 23.670 22.860 25.090 23.030 ;
        RECT 25.900 22.860 26.320 23.070 ;
        RECT 26.830 22.860 27.250 23.070 ;
        RECT 22.730 22.420 24.310 22.590 ;
        RECT 25.520 22.470 25.690 22.800 ;
        RECT 19.560 21.650 19.730 21.980 ;
        RECT 20.970 21.860 22.550 22.030 ;
        RECT 18.030 21.380 18.450 21.590 ;
        RECT 18.920 21.380 19.340 21.590 ;
        RECT 20.150 21.420 21.610 21.590 ;
        RECT 18.100 21.320 18.360 21.380 ;
        RECT 19.010 21.320 19.270 21.380 ;
        RECT 20.610 21.360 20.900 21.420 ;
        RECT 22.130 21.250 22.550 21.590 ;
        RECT 22.810 21.550 22.980 22.420 ;
        RECT 23.360 21.550 23.530 22.240 ;
        RECT 27.500 22.200 27.670 22.890 ;
        RECT 28.040 22.030 28.210 22.900 ;
        RECT 28.480 22.860 28.900 23.140 ;
        RECT 30.120 23.030 30.290 23.360 ;
        RECT 31.740 23.070 32.000 23.160 ;
        RECT 32.650 23.070 32.910 23.160 ;
        RECT 29.420 22.860 30.840 23.030 ;
        RECT 31.650 22.860 32.070 23.070 ;
        RECT 32.580 22.860 33.000 23.070 ;
        RECT 28.480 22.420 30.060 22.590 ;
        RECT 31.270 22.470 31.440 22.800 ;
        RECT 25.310 21.650 25.480 21.980 ;
        RECT 26.720 21.860 28.300 22.030 ;
        RECT 23.780 21.380 24.200 21.590 ;
        RECT 24.670 21.380 25.090 21.590 ;
        RECT 25.900 21.420 27.360 21.590 ;
        RECT 23.850 21.320 24.110 21.380 ;
        RECT 24.760 21.320 25.020 21.380 ;
        RECT 26.360 21.360 26.650 21.420 ;
        RECT 27.880 21.250 28.300 21.590 ;
        RECT 28.560 21.550 28.730 22.420 ;
        RECT 29.110 21.550 29.280 22.240 ;
        RECT 33.250 22.200 33.420 22.890 ;
        RECT 33.790 22.030 33.960 22.900 ;
        RECT 34.230 22.860 34.650 23.140 ;
        RECT 35.870 23.030 36.040 23.360 ;
        RECT 37.490 23.070 37.750 23.160 ;
        RECT 38.400 23.070 38.660 23.160 ;
        RECT 35.170 22.860 36.590 23.030 ;
        RECT 37.400 22.860 37.820 23.070 ;
        RECT 38.330 22.860 38.750 23.070 ;
        RECT 34.230 22.420 35.810 22.590 ;
        RECT 37.020 22.470 37.190 22.800 ;
        RECT 31.060 21.650 31.230 21.980 ;
        RECT 32.470 21.860 34.050 22.030 ;
        RECT 29.530 21.380 29.950 21.590 ;
        RECT 30.420 21.380 30.840 21.590 ;
        RECT 31.650 21.420 33.110 21.590 ;
        RECT 29.600 21.320 29.860 21.380 ;
        RECT 30.510 21.320 30.770 21.380 ;
        RECT 32.110 21.360 32.400 21.420 ;
        RECT 33.630 21.250 34.050 21.590 ;
        RECT 34.310 21.550 34.480 22.420 ;
        RECT 34.860 21.550 35.030 22.240 ;
        RECT 39.000 22.200 39.170 22.890 ;
        RECT 39.540 22.030 39.710 22.900 ;
        RECT 39.980 22.860 40.400 23.140 ;
        RECT 41.620 23.030 41.790 23.360 ;
        RECT 43.240 23.070 43.500 23.160 ;
        RECT 44.150 23.070 44.410 23.160 ;
        RECT 40.920 22.860 42.340 23.030 ;
        RECT 43.150 22.860 43.570 23.070 ;
        RECT 44.080 22.860 44.500 23.070 ;
        RECT 39.980 22.420 41.560 22.590 ;
        RECT 42.770 22.470 42.940 22.800 ;
        RECT 36.810 21.650 36.980 21.980 ;
        RECT 38.220 21.860 39.800 22.030 ;
        RECT 35.280 21.380 35.700 21.590 ;
        RECT 36.170 21.380 36.590 21.590 ;
        RECT 37.400 21.420 38.860 21.590 ;
        RECT 35.350 21.320 35.610 21.380 ;
        RECT 36.260 21.320 36.520 21.380 ;
        RECT 37.860 21.360 38.150 21.420 ;
        RECT 39.380 21.250 39.800 21.590 ;
        RECT 40.060 21.550 40.230 22.420 ;
        RECT 40.610 21.550 40.780 22.240 ;
        RECT 44.750 22.200 44.920 22.890 ;
        RECT 45.290 22.030 45.460 22.900 ;
        RECT 45.730 22.860 46.150 23.140 ;
        RECT 47.370 23.030 47.540 23.360 ;
        RECT 48.990 23.070 49.250 23.160 ;
        RECT 49.900 23.070 50.160 23.160 ;
        RECT 46.670 22.860 48.090 23.030 ;
        RECT 48.900 22.860 49.320 23.070 ;
        RECT 49.830 22.860 50.250 23.070 ;
        RECT 45.730 22.420 47.310 22.590 ;
        RECT 48.520 22.470 48.690 22.800 ;
        RECT 42.560 21.650 42.730 21.980 ;
        RECT 43.970 21.860 45.550 22.030 ;
        RECT 41.030 21.380 41.450 21.590 ;
        RECT 41.920 21.380 42.340 21.590 ;
        RECT 43.150 21.420 44.610 21.590 ;
        RECT 41.100 21.320 41.360 21.380 ;
        RECT 42.010 21.320 42.270 21.380 ;
        RECT 43.610 21.360 43.900 21.420 ;
        RECT 45.130 21.250 45.550 21.590 ;
        RECT 45.810 21.550 45.980 22.420 ;
        RECT 46.360 21.550 46.530 22.240 ;
        RECT 50.500 22.200 50.670 22.890 ;
        RECT 51.040 22.030 51.210 22.900 ;
        RECT 51.480 22.860 51.900 23.140 ;
        RECT 53.120 23.030 53.290 23.360 ;
        RECT 54.740 23.070 55.000 23.160 ;
        RECT 55.650 23.070 55.910 23.160 ;
        RECT 52.420 22.860 53.840 23.030 ;
        RECT 54.650 22.860 55.070 23.070 ;
        RECT 55.580 22.860 56.000 23.070 ;
        RECT 51.480 22.420 53.060 22.590 ;
        RECT 54.270 22.470 54.440 22.800 ;
        RECT 48.310 21.650 48.480 21.980 ;
        RECT 49.720 21.860 51.300 22.030 ;
        RECT 46.780 21.380 47.200 21.590 ;
        RECT 47.670 21.380 48.090 21.590 ;
        RECT 48.900 21.420 50.360 21.590 ;
        RECT 46.850 21.320 47.110 21.380 ;
        RECT 47.760 21.320 48.020 21.380 ;
        RECT 49.360 21.360 49.650 21.420 ;
        RECT 50.880 21.250 51.300 21.590 ;
        RECT 51.560 21.550 51.730 22.420 ;
        RECT 52.110 21.550 52.280 22.240 ;
        RECT 56.250 22.200 56.420 22.890 ;
        RECT 56.790 22.030 56.960 22.900 ;
        RECT 57.230 22.860 57.650 23.140 ;
        RECT 58.870 23.030 59.040 23.360 ;
        RECT 60.490 23.070 60.750 23.160 ;
        RECT 61.400 23.070 61.660 23.160 ;
        RECT 58.170 22.860 59.590 23.030 ;
        RECT 60.400 22.860 60.820 23.070 ;
        RECT 61.330 22.860 61.750 23.070 ;
        RECT 57.230 22.420 58.810 22.590 ;
        RECT 60.020 22.470 60.190 22.800 ;
        RECT 54.060 21.650 54.230 21.980 ;
        RECT 55.470 21.860 57.050 22.030 ;
        RECT 52.530 21.380 52.950 21.590 ;
        RECT 53.420 21.380 53.840 21.590 ;
        RECT 54.650 21.420 56.110 21.590 ;
        RECT 52.600 21.320 52.860 21.380 ;
        RECT 53.510 21.320 53.770 21.380 ;
        RECT 55.110 21.360 55.400 21.420 ;
        RECT 56.630 21.250 57.050 21.590 ;
        RECT 57.310 21.550 57.480 22.420 ;
        RECT 57.860 21.550 58.030 22.240 ;
        RECT 62.000 22.200 62.170 22.890 ;
        RECT 62.540 22.030 62.710 22.900 ;
        RECT 62.980 22.860 63.400 23.140 ;
        RECT 64.620 23.030 64.790 23.360 ;
        RECT 66.240 23.070 66.500 23.160 ;
        RECT 67.150 23.070 67.410 23.160 ;
        RECT 63.920 22.860 65.340 23.030 ;
        RECT 66.150 22.860 66.570 23.070 ;
        RECT 67.080 22.860 67.500 23.070 ;
        RECT 62.980 22.420 64.560 22.590 ;
        RECT 65.770 22.470 65.940 22.800 ;
        RECT 59.810 21.650 59.980 21.980 ;
        RECT 61.220 21.860 62.800 22.030 ;
        RECT 58.280 21.380 58.700 21.590 ;
        RECT 59.170 21.380 59.590 21.590 ;
        RECT 60.400 21.420 61.860 21.590 ;
        RECT 58.350 21.320 58.610 21.380 ;
        RECT 59.260 21.320 59.520 21.380 ;
        RECT 60.860 21.360 61.150 21.420 ;
        RECT 62.380 21.250 62.800 21.590 ;
        RECT 63.060 21.550 63.230 22.420 ;
        RECT 63.610 21.550 63.780 22.240 ;
        RECT 67.750 22.200 67.920 22.890 ;
        RECT 68.290 22.030 68.460 22.900 ;
        RECT 68.730 22.860 69.150 23.140 ;
        RECT 70.370 23.030 70.540 23.360 ;
        RECT 71.990 23.070 72.250 23.160 ;
        RECT 72.900 23.070 73.160 23.160 ;
        RECT 69.670 22.860 71.090 23.030 ;
        RECT 71.900 22.860 72.320 23.070 ;
        RECT 72.830 22.860 73.250 23.070 ;
        RECT 68.730 22.420 70.310 22.590 ;
        RECT 71.520 22.470 71.690 22.800 ;
        RECT 65.560 21.650 65.730 21.980 ;
        RECT 66.970 21.860 68.550 22.030 ;
        RECT 64.030 21.380 64.450 21.590 ;
        RECT 64.920 21.380 65.340 21.590 ;
        RECT 66.150 21.420 67.610 21.590 ;
        RECT 64.100 21.320 64.360 21.380 ;
        RECT 65.010 21.320 65.270 21.380 ;
        RECT 66.610 21.360 66.900 21.420 ;
        RECT 68.130 21.250 68.550 21.590 ;
        RECT 68.810 21.550 68.980 22.420 ;
        RECT 69.360 21.550 69.530 22.240 ;
        RECT 73.500 22.200 73.670 22.890 ;
        RECT 74.040 22.030 74.210 22.900 ;
        RECT 74.480 22.860 74.900 23.140 ;
        RECT 76.120 23.030 76.290 23.360 ;
        RECT 77.740 23.070 78.000 23.160 ;
        RECT 78.650 23.070 78.910 23.160 ;
        RECT 75.420 22.860 76.840 23.030 ;
        RECT 77.650 22.860 78.070 23.070 ;
        RECT 78.580 22.860 79.000 23.070 ;
        RECT 74.480 22.420 76.060 22.590 ;
        RECT 77.270 22.470 77.440 22.800 ;
        RECT 71.310 21.650 71.480 21.980 ;
        RECT 72.720 21.860 74.300 22.030 ;
        RECT 69.780 21.380 70.200 21.590 ;
        RECT 70.670 21.380 71.090 21.590 ;
        RECT 71.900 21.420 73.360 21.590 ;
        RECT 69.850 21.320 70.110 21.380 ;
        RECT 70.760 21.320 71.020 21.380 ;
        RECT 72.360 21.360 72.650 21.420 ;
        RECT 73.880 21.250 74.300 21.590 ;
        RECT 74.560 21.550 74.730 22.420 ;
        RECT 75.110 21.550 75.280 22.240 ;
        RECT 79.250 22.200 79.420 22.890 ;
        RECT 79.790 22.030 79.960 22.900 ;
        RECT 80.230 22.860 80.650 23.140 ;
        RECT 81.870 23.030 82.040 23.360 ;
        RECT 83.490 23.070 83.750 23.160 ;
        RECT 84.400 23.070 84.660 23.160 ;
        RECT 81.170 22.860 82.590 23.030 ;
        RECT 83.400 22.860 83.820 23.070 ;
        RECT 84.330 22.860 84.750 23.070 ;
        RECT 80.230 22.420 81.810 22.590 ;
        RECT 83.020 22.470 83.190 22.800 ;
        RECT 77.060 21.650 77.230 21.980 ;
        RECT 78.470 21.860 80.050 22.030 ;
        RECT 75.530 21.380 75.950 21.590 ;
        RECT 76.420 21.380 76.840 21.590 ;
        RECT 77.650 21.420 79.110 21.590 ;
        RECT 75.600 21.320 75.860 21.380 ;
        RECT 76.510 21.320 76.770 21.380 ;
        RECT 78.110 21.360 78.400 21.420 ;
        RECT 79.630 21.250 80.050 21.590 ;
        RECT 80.310 21.550 80.480 22.420 ;
        RECT 80.860 21.550 81.030 22.240 ;
        RECT 85.000 22.200 85.170 22.890 ;
        RECT 85.540 22.030 85.710 22.900 ;
        RECT 85.980 22.860 86.400 23.140 ;
        RECT 87.620 23.030 87.790 23.360 ;
        RECT 89.240 23.070 89.500 23.160 ;
        RECT 90.150 23.070 90.410 23.160 ;
        RECT 86.920 22.860 88.340 23.030 ;
        RECT 89.150 22.860 89.570 23.070 ;
        RECT 90.080 22.860 90.500 23.070 ;
        RECT 85.980 22.420 87.560 22.590 ;
        RECT 88.770 22.470 88.940 22.800 ;
        RECT 82.810 21.650 82.980 21.980 ;
        RECT 84.220 21.860 85.800 22.030 ;
        RECT 81.280 21.380 81.700 21.590 ;
        RECT 82.170 21.380 82.590 21.590 ;
        RECT 83.400 21.420 84.860 21.590 ;
        RECT 81.350 21.320 81.610 21.380 ;
        RECT 82.260 21.320 82.520 21.380 ;
        RECT 83.860 21.360 84.150 21.420 ;
        RECT 85.380 21.250 85.800 21.590 ;
        RECT 86.060 21.550 86.230 22.420 ;
        RECT 86.610 21.550 86.780 22.240 ;
        RECT 90.750 22.200 90.920 22.890 ;
        RECT 91.290 22.030 91.460 22.900 ;
        RECT 91.730 22.860 92.150 23.140 ;
        RECT 93.370 23.030 93.540 23.360 ;
        RECT 92.670 22.860 94.090 23.030 ;
        RECT 91.730 22.420 93.310 22.590 ;
        RECT 88.560 21.650 88.730 21.980 ;
        RECT 89.970 21.860 91.550 22.030 ;
        RECT 87.030 21.380 87.450 21.590 ;
        RECT 87.920 21.380 88.340 21.590 ;
        RECT 89.150 21.420 90.610 21.590 ;
        RECT 87.100 21.320 87.360 21.380 ;
        RECT 88.010 21.320 88.270 21.380 ;
        RECT 89.610 21.360 89.900 21.420 ;
        RECT 91.130 21.250 91.550 21.590 ;
        RECT 91.810 21.550 91.980 22.420 ;
        RECT 92.360 21.550 92.530 22.240 ;
        RECT 94.310 21.650 94.480 21.980 ;
        RECT 92.780 21.380 93.200 21.590 ;
        RECT 93.670 21.380 94.090 21.590 ;
        RECT 92.850 21.320 93.110 21.380 ;
        RECT 93.760 21.320 94.020 21.380 ;
        RECT 2.990 20.660 3.250 20.750 ;
        RECT 3.900 20.660 4.160 20.750 ;
        RECT 2.900 20.450 3.320 20.660 ;
        RECT 3.830 20.450 4.250 20.660 ;
        RECT 2.520 20.060 2.690 20.390 ;
        RECT 4.500 19.790 4.670 20.480 ;
        RECT 5.040 19.620 5.210 20.490 ;
        RECT 5.480 20.450 5.900 20.730 ;
        RECT 7.120 20.620 7.290 20.950 ;
        RECT 8.740 20.660 9.000 20.750 ;
        RECT 9.650 20.660 9.910 20.750 ;
        RECT 6.420 20.450 7.840 20.620 ;
        RECT 8.650 20.450 9.070 20.660 ;
        RECT 9.580 20.450 10.000 20.660 ;
        RECT 5.480 20.010 7.060 20.180 ;
        RECT 8.270 20.060 8.440 20.390 ;
        RECT 3.720 19.450 5.300 19.620 ;
        RECT 2.900 19.010 4.360 19.180 ;
        RECT 3.360 18.950 3.650 19.010 ;
        RECT 4.880 18.840 5.300 19.180 ;
        RECT 5.560 19.140 5.730 20.010 ;
        RECT 6.110 19.140 6.280 19.830 ;
        RECT 10.250 19.790 10.420 20.480 ;
        RECT 10.790 19.620 10.960 20.490 ;
        RECT 11.230 20.450 11.650 20.730 ;
        RECT 12.870 20.620 13.040 20.950 ;
        RECT 14.490 20.660 14.750 20.750 ;
        RECT 15.400 20.660 15.660 20.750 ;
        RECT 12.170 20.450 13.590 20.620 ;
        RECT 14.400 20.450 14.820 20.660 ;
        RECT 15.330 20.450 15.750 20.660 ;
        RECT 11.230 20.010 12.810 20.180 ;
        RECT 14.020 20.060 14.190 20.390 ;
        RECT 8.060 19.240 8.230 19.570 ;
        RECT 9.470 19.450 11.050 19.620 ;
        RECT 6.530 18.970 6.950 19.180 ;
        RECT 7.420 18.970 7.840 19.180 ;
        RECT 8.650 19.010 10.110 19.180 ;
        RECT 6.600 18.910 6.860 18.970 ;
        RECT 7.510 18.910 7.770 18.970 ;
        RECT 9.110 18.950 9.400 19.010 ;
        RECT 10.630 18.840 11.050 19.180 ;
        RECT 11.310 19.140 11.480 20.010 ;
        RECT 11.860 19.140 12.030 19.830 ;
        RECT 16.000 19.790 16.170 20.480 ;
        RECT 16.540 19.620 16.710 20.490 ;
        RECT 16.980 20.450 17.400 20.730 ;
        RECT 18.620 20.620 18.790 20.950 ;
        RECT 20.240 20.660 20.500 20.750 ;
        RECT 21.150 20.660 21.410 20.750 ;
        RECT 17.920 20.450 19.340 20.620 ;
        RECT 20.150 20.450 20.570 20.660 ;
        RECT 21.080 20.450 21.500 20.660 ;
        RECT 16.980 20.010 18.560 20.180 ;
        RECT 19.770 20.060 19.940 20.390 ;
        RECT 13.810 19.240 13.980 19.570 ;
        RECT 15.220 19.450 16.800 19.620 ;
        RECT 12.280 18.970 12.700 19.180 ;
        RECT 13.170 18.970 13.590 19.180 ;
        RECT 14.400 19.010 15.860 19.180 ;
        RECT 12.350 18.910 12.610 18.970 ;
        RECT 13.260 18.910 13.520 18.970 ;
        RECT 14.860 18.950 15.150 19.010 ;
        RECT 16.380 18.840 16.800 19.180 ;
        RECT 17.060 19.140 17.230 20.010 ;
        RECT 17.610 19.140 17.780 19.830 ;
        RECT 21.750 19.790 21.920 20.480 ;
        RECT 22.290 19.620 22.460 20.490 ;
        RECT 22.730 20.450 23.150 20.730 ;
        RECT 24.370 20.620 24.540 20.950 ;
        RECT 25.990 20.660 26.250 20.750 ;
        RECT 26.900 20.660 27.160 20.750 ;
        RECT 23.670 20.450 25.090 20.620 ;
        RECT 25.900 20.450 26.320 20.660 ;
        RECT 26.830 20.450 27.250 20.660 ;
        RECT 22.730 20.010 24.310 20.180 ;
        RECT 25.520 20.060 25.690 20.390 ;
        RECT 19.560 19.240 19.730 19.570 ;
        RECT 20.970 19.450 22.550 19.620 ;
        RECT 18.030 18.970 18.450 19.180 ;
        RECT 18.920 18.970 19.340 19.180 ;
        RECT 20.150 19.010 21.610 19.180 ;
        RECT 18.100 18.910 18.360 18.970 ;
        RECT 19.010 18.910 19.270 18.970 ;
        RECT 20.610 18.950 20.900 19.010 ;
        RECT 22.130 18.840 22.550 19.180 ;
        RECT 22.810 19.140 22.980 20.010 ;
        RECT 23.360 19.140 23.530 19.830 ;
        RECT 27.500 19.790 27.670 20.480 ;
        RECT 28.040 19.620 28.210 20.490 ;
        RECT 28.480 20.450 28.900 20.730 ;
        RECT 30.120 20.620 30.290 20.950 ;
        RECT 31.740 20.660 32.000 20.750 ;
        RECT 32.650 20.660 32.910 20.750 ;
        RECT 29.420 20.450 30.840 20.620 ;
        RECT 31.650 20.450 32.070 20.660 ;
        RECT 32.580 20.450 33.000 20.660 ;
        RECT 28.480 20.010 30.060 20.180 ;
        RECT 31.270 20.060 31.440 20.390 ;
        RECT 25.310 19.240 25.480 19.570 ;
        RECT 26.720 19.450 28.300 19.620 ;
        RECT 23.780 18.970 24.200 19.180 ;
        RECT 24.670 18.970 25.090 19.180 ;
        RECT 25.900 19.010 27.360 19.180 ;
        RECT 23.850 18.910 24.110 18.970 ;
        RECT 24.760 18.910 25.020 18.970 ;
        RECT 26.360 18.950 26.650 19.010 ;
        RECT 27.880 18.840 28.300 19.180 ;
        RECT 28.560 19.140 28.730 20.010 ;
        RECT 29.110 19.140 29.280 19.830 ;
        RECT 33.250 19.790 33.420 20.480 ;
        RECT 33.790 19.620 33.960 20.490 ;
        RECT 34.230 20.450 34.650 20.730 ;
        RECT 35.870 20.620 36.040 20.950 ;
        RECT 37.490 20.660 37.750 20.750 ;
        RECT 38.400 20.660 38.660 20.750 ;
        RECT 35.170 20.450 36.590 20.620 ;
        RECT 37.400 20.450 37.820 20.660 ;
        RECT 38.330 20.450 38.750 20.660 ;
        RECT 34.230 20.010 35.810 20.180 ;
        RECT 37.020 20.060 37.190 20.390 ;
        RECT 31.060 19.240 31.230 19.570 ;
        RECT 32.470 19.450 34.050 19.620 ;
        RECT 29.530 18.970 29.950 19.180 ;
        RECT 30.420 18.970 30.840 19.180 ;
        RECT 31.650 19.010 33.110 19.180 ;
        RECT 29.600 18.910 29.860 18.970 ;
        RECT 30.510 18.910 30.770 18.970 ;
        RECT 32.110 18.950 32.400 19.010 ;
        RECT 33.630 18.840 34.050 19.180 ;
        RECT 34.310 19.140 34.480 20.010 ;
        RECT 34.860 19.140 35.030 19.830 ;
        RECT 39.000 19.790 39.170 20.480 ;
        RECT 39.540 19.620 39.710 20.490 ;
        RECT 39.980 20.450 40.400 20.730 ;
        RECT 41.620 20.620 41.790 20.950 ;
        RECT 43.240 20.660 43.500 20.750 ;
        RECT 44.150 20.660 44.410 20.750 ;
        RECT 40.920 20.450 42.340 20.620 ;
        RECT 43.150 20.450 43.570 20.660 ;
        RECT 44.080 20.450 44.500 20.660 ;
        RECT 39.980 20.010 41.560 20.180 ;
        RECT 42.770 20.060 42.940 20.390 ;
        RECT 36.810 19.240 36.980 19.570 ;
        RECT 38.220 19.450 39.800 19.620 ;
        RECT 35.280 18.970 35.700 19.180 ;
        RECT 36.170 18.970 36.590 19.180 ;
        RECT 37.400 19.010 38.860 19.180 ;
        RECT 35.350 18.910 35.610 18.970 ;
        RECT 36.260 18.910 36.520 18.970 ;
        RECT 37.860 18.950 38.150 19.010 ;
        RECT 39.380 18.840 39.800 19.180 ;
        RECT 40.060 19.140 40.230 20.010 ;
        RECT 40.610 19.140 40.780 19.830 ;
        RECT 44.750 19.790 44.920 20.480 ;
        RECT 45.290 19.620 45.460 20.490 ;
        RECT 45.730 20.450 46.150 20.730 ;
        RECT 47.370 20.620 47.540 20.950 ;
        RECT 48.990 20.660 49.250 20.750 ;
        RECT 49.900 20.660 50.160 20.750 ;
        RECT 46.670 20.450 48.090 20.620 ;
        RECT 48.900 20.450 49.320 20.660 ;
        RECT 49.830 20.450 50.250 20.660 ;
        RECT 45.730 20.010 47.310 20.180 ;
        RECT 48.520 20.060 48.690 20.390 ;
        RECT 42.560 19.240 42.730 19.570 ;
        RECT 43.970 19.450 45.550 19.620 ;
        RECT 41.030 18.970 41.450 19.180 ;
        RECT 41.920 18.970 42.340 19.180 ;
        RECT 43.150 19.010 44.610 19.180 ;
        RECT 41.100 18.910 41.360 18.970 ;
        RECT 42.010 18.910 42.270 18.970 ;
        RECT 43.610 18.950 43.900 19.010 ;
        RECT 45.130 18.840 45.550 19.180 ;
        RECT 45.810 19.140 45.980 20.010 ;
        RECT 46.360 19.140 46.530 19.830 ;
        RECT 50.500 19.790 50.670 20.480 ;
        RECT 51.040 19.620 51.210 20.490 ;
        RECT 51.480 20.450 51.900 20.730 ;
        RECT 53.120 20.620 53.290 20.950 ;
        RECT 54.740 20.660 55.000 20.750 ;
        RECT 55.650 20.660 55.910 20.750 ;
        RECT 52.420 20.450 53.840 20.620 ;
        RECT 54.650 20.450 55.070 20.660 ;
        RECT 55.580 20.450 56.000 20.660 ;
        RECT 51.480 20.010 53.060 20.180 ;
        RECT 54.270 20.060 54.440 20.390 ;
        RECT 48.310 19.240 48.480 19.570 ;
        RECT 49.720 19.450 51.300 19.620 ;
        RECT 46.780 18.970 47.200 19.180 ;
        RECT 47.670 18.970 48.090 19.180 ;
        RECT 48.900 19.010 50.360 19.180 ;
        RECT 46.850 18.910 47.110 18.970 ;
        RECT 47.760 18.910 48.020 18.970 ;
        RECT 49.360 18.950 49.650 19.010 ;
        RECT 50.880 18.840 51.300 19.180 ;
        RECT 51.560 19.140 51.730 20.010 ;
        RECT 52.110 19.140 52.280 19.830 ;
        RECT 56.250 19.790 56.420 20.480 ;
        RECT 56.790 19.620 56.960 20.490 ;
        RECT 57.230 20.450 57.650 20.730 ;
        RECT 58.870 20.620 59.040 20.950 ;
        RECT 60.490 20.660 60.750 20.750 ;
        RECT 61.400 20.660 61.660 20.750 ;
        RECT 58.170 20.450 59.590 20.620 ;
        RECT 60.400 20.450 60.820 20.660 ;
        RECT 61.330 20.450 61.750 20.660 ;
        RECT 57.230 20.010 58.810 20.180 ;
        RECT 60.020 20.060 60.190 20.390 ;
        RECT 54.060 19.240 54.230 19.570 ;
        RECT 55.470 19.450 57.050 19.620 ;
        RECT 52.530 18.970 52.950 19.180 ;
        RECT 53.420 18.970 53.840 19.180 ;
        RECT 54.650 19.010 56.110 19.180 ;
        RECT 52.600 18.910 52.860 18.970 ;
        RECT 53.510 18.910 53.770 18.970 ;
        RECT 55.110 18.950 55.400 19.010 ;
        RECT 56.630 18.840 57.050 19.180 ;
        RECT 57.310 19.140 57.480 20.010 ;
        RECT 57.860 19.140 58.030 19.830 ;
        RECT 62.000 19.790 62.170 20.480 ;
        RECT 62.540 19.620 62.710 20.490 ;
        RECT 62.980 20.450 63.400 20.730 ;
        RECT 64.620 20.620 64.790 20.950 ;
        RECT 66.240 20.660 66.500 20.750 ;
        RECT 67.150 20.660 67.410 20.750 ;
        RECT 63.920 20.450 65.340 20.620 ;
        RECT 66.150 20.450 66.570 20.660 ;
        RECT 67.080 20.450 67.500 20.660 ;
        RECT 62.980 20.010 64.560 20.180 ;
        RECT 65.770 20.060 65.940 20.390 ;
        RECT 59.810 19.240 59.980 19.570 ;
        RECT 61.220 19.450 62.800 19.620 ;
        RECT 58.280 18.970 58.700 19.180 ;
        RECT 59.170 18.970 59.590 19.180 ;
        RECT 60.400 19.010 61.860 19.180 ;
        RECT 58.350 18.910 58.610 18.970 ;
        RECT 59.260 18.910 59.520 18.970 ;
        RECT 60.860 18.950 61.150 19.010 ;
        RECT 62.380 18.840 62.800 19.180 ;
        RECT 63.060 19.140 63.230 20.010 ;
        RECT 63.610 19.140 63.780 19.830 ;
        RECT 67.750 19.790 67.920 20.480 ;
        RECT 68.290 19.620 68.460 20.490 ;
        RECT 68.730 20.450 69.150 20.730 ;
        RECT 70.370 20.620 70.540 20.950 ;
        RECT 71.990 20.660 72.250 20.750 ;
        RECT 72.900 20.660 73.160 20.750 ;
        RECT 69.670 20.450 71.090 20.620 ;
        RECT 71.900 20.450 72.320 20.660 ;
        RECT 72.830 20.450 73.250 20.660 ;
        RECT 68.730 20.010 70.310 20.180 ;
        RECT 71.520 20.060 71.690 20.390 ;
        RECT 65.560 19.240 65.730 19.570 ;
        RECT 66.970 19.450 68.550 19.620 ;
        RECT 64.030 18.970 64.450 19.180 ;
        RECT 64.920 18.970 65.340 19.180 ;
        RECT 66.150 19.010 67.610 19.180 ;
        RECT 64.100 18.910 64.360 18.970 ;
        RECT 65.010 18.910 65.270 18.970 ;
        RECT 66.610 18.950 66.900 19.010 ;
        RECT 68.130 18.840 68.550 19.180 ;
        RECT 68.810 19.140 68.980 20.010 ;
        RECT 69.360 19.140 69.530 19.830 ;
        RECT 73.500 19.790 73.670 20.480 ;
        RECT 74.040 19.620 74.210 20.490 ;
        RECT 74.480 20.450 74.900 20.730 ;
        RECT 76.120 20.620 76.290 20.950 ;
        RECT 77.740 20.660 78.000 20.750 ;
        RECT 78.650 20.660 78.910 20.750 ;
        RECT 75.420 20.450 76.840 20.620 ;
        RECT 77.650 20.450 78.070 20.660 ;
        RECT 78.580 20.450 79.000 20.660 ;
        RECT 74.480 20.010 76.060 20.180 ;
        RECT 77.270 20.060 77.440 20.390 ;
        RECT 71.310 19.240 71.480 19.570 ;
        RECT 72.720 19.450 74.300 19.620 ;
        RECT 69.780 18.970 70.200 19.180 ;
        RECT 70.670 18.970 71.090 19.180 ;
        RECT 71.900 19.010 73.360 19.180 ;
        RECT 69.850 18.910 70.110 18.970 ;
        RECT 70.760 18.910 71.020 18.970 ;
        RECT 72.360 18.950 72.650 19.010 ;
        RECT 73.880 18.840 74.300 19.180 ;
        RECT 74.560 19.140 74.730 20.010 ;
        RECT 75.110 19.140 75.280 19.830 ;
        RECT 79.250 19.790 79.420 20.480 ;
        RECT 79.790 19.620 79.960 20.490 ;
        RECT 80.230 20.450 80.650 20.730 ;
        RECT 81.870 20.620 82.040 20.950 ;
        RECT 83.490 20.660 83.750 20.750 ;
        RECT 84.400 20.660 84.660 20.750 ;
        RECT 81.170 20.450 82.590 20.620 ;
        RECT 83.400 20.450 83.820 20.660 ;
        RECT 84.330 20.450 84.750 20.660 ;
        RECT 80.230 20.010 81.810 20.180 ;
        RECT 83.020 20.060 83.190 20.390 ;
        RECT 77.060 19.240 77.230 19.570 ;
        RECT 78.470 19.450 80.050 19.620 ;
        RECT 75.530 18.970 75.950 19.180 ;
        RECT 76.420 18.970 76.840 19.180 ;
        RECT 77.650 19.010 79.110 19.180 ;
        RECT 75.600 18.910 75.860 18.970 ;
        RECT 76.510 18.910 76.770 18.970 ;
        RECT 78.110 18.950 78.400 19.010 ;
        RECT 79.630 18.840 80.050 19.180 ;
        RECT 80.310 19.140 80.480 20.010 ;
        RECT 80.860 19.140 81.030 19.830 ;
        RECT 85.000 19.790 85.170 20.480 ;
        RECT 85.540 19.620 85.710 20.490 ;
        RECT 85.980 20.450 86.400 20.730 ;
        RECT 87.620 20.620 87.790 20.950 ;
        RECT 89.240 20.660 89.500 20.750 ;
        RECT 90.150 20.660 90.410 20.750 ;
        RECT 86.920 20.450 88.340 20.620 ;
        RECT 89.150 20.450 89.570 20.660 ;
        RECT 90.080 20.450 90.500 20.660 ;
        RECT 85.980 20.010 87.560 20.180 ;
        RECT 88.770 20.060 88.940 20.390 ;
        RECT 82.810 19.240 82.980 19.570 ;
        RECT 84.220 19.450 85.800 19.620 ;
        RECT 81.280 18.970 81.700 19.180 ;
        RECT 82.170 18.970 82.590 19.180 ;
        RECT 83.400 19.010 84.860 19.180 ;
        RECT 81.350 18.910 81.610 18.970 ;
        RECT 82.260 18.910 82.520 18.970 ;
        RECT 83.860 18.950 84.150 19.010 ;
        RECT 85.380 18.840 85.800 19.180 ;
        RECT 86.060 19.140 86.230 20.010 ;
        RECT 86.610 19.140 86.780 19.830 ;
        RECT 90.750 19.790 90.920 20.480 ;
        RECT 91.290 19.620 91.460 20.490 ;
        RECT 91.730 20.450 92.150 20.730 ;
        RECT 93.370 20.620 93.540 20.950 ;
        RECT 92.670 20.450 94.090 20.620 ;
        RECT 91.730 20.010 93.310 20.180 ;
        RECT 88.560 19.240 88.730 19.570 ;
        RECT 89.970 19.450 91.550 19.620 ;
        RECT 87.030 18.970 87.450 19.180 ;
        RECT 87.920 18.970 88.340 19.180 ;
        RECT 89.150 19.010 90.610 19.180 ;
        RECT 87.100 18.910 87.360 18.970 ;
        RECT 88.010 18.910 88.270 18.970 ;
        RECT 89.610 18.950 89.900 19.010 ;
        RECT 91.130 18.840 91.550 19.180 ;
        RECT 91.810 19.140 91.980 20.010 ;
        RECT 92.360 19.140 92.530 19.830 ;
        RECT 94.310 19.240 94.480 19.570 ;
        RECT 92.780 18.970 93.200 19.180 ;
        RECT 93.670 18.970 94.090 19.180 ;
        RECT 92.850 18.910 93.110 18.970 ;
        RECT 93.760 18.910 94.020 18.970 ;
        RECT 2.990 18.250 3.250 18.340 ;
        RECT 3.900 18.250 4.160 18.340 ;
        RECT 2.900 18.040 3.320 18.250 ;
        RECT 3.830 18.040 4.250 18.250 ;
        RECT 2.520 17.650 2.690 17.980 ;
        RECT 4.500 17.380 4.670 18.070 ;
        RECT 5.040 17.210 5.210 18.080 ;
        RECT 5.480 18.040 5.900 18.320 ;
        RECT 7.120 18.210 7.290 18.540 ;
        RECT 8.740 18.250 9.000 18.340 ;
        RECT 9.650 18.250 9.910 18.340 ;
        RECT 6.420 18.040 7.840 18.210 ;
        RECT 8.650 18.040 9.070 18.250 ;
        RECT 9.580 18.040 10.000 18.250 ;
        RECT 5.480 17.600 7.060 17.770 ;
        RECT 8.270 17.650 8.440 17.980 ;
        RECT 3.720 17.040 5.300 17.210 ;
        RECT 2.900 16.600 4.360 16.770 ;
        RECT 3.360 16.540 3.650 16.600 ;
        RECT 4.880 16.430 5.300 16.770 ;
        RECT 5.560 16.730 5.730 17.600 ;
        RECT 6.110 16.730 6.280 17.420 ;
        RECT 10.250 17.380 10.420 18.070 ;
        RECT 10.790 17.210 10.960 18.080 ;
        RECT 11.230 18.040 11.650 18.320 ;
        RECT 12.870 18.210 13.040 18.540 ;
        RECT 14.490 18.250 14.750 18.340 ;
        RECT 15.400 18.250 15.660 18.340 ;
        RECT 12.170 18.040 13.590 18.210 ;
        RECT 14.400 18.040 14.820 18.250 ;
        RECT 15.330 18.040 15.750 18.250 ;
        RECT 11.230 17.600 12.810 17.770 ;
        RECT 14.020 17.650 14.190 17.980 ;
        RECT 8.060 16.830 8.230 17.160 ;
        RECT 9.470 17.040 11.050 17.210 ;
        RECT 6.530 16.560 6.950 16.770 ;
        RECT 7.420 16.560 7.840 16.770 ;
        RECT 8.650 16.600 10.110 16.770 ;
        RECT 6.600 16.500 6.860 16.560 ;
        RECT 7.510 16.500 7.770 16.560 ;
        RECT 9.110 16.540 9.400 16.600 ;
        RECT 10.630 16.430 11.050 16.770 ;
        RECT 11.310 16.730 11.480 17.600 ;
        RECT 11.860 16.730 12.030 17.420 ;
        RECT 16.000 17.380 16.170 18.070 ;
        RECT 16.540 17.210 16.710 18.080 ;
        RECT 16.980 18.040 17.400 18.320 ;
        RECT 18.620 18.210 18.790 18.540 ;
        RECT 20.240 18.250 20.500 18.340 ;
        RECT 21.150 18.250 21.410 18.340 ;
        RECT 17.920 18.040 19.340 18.210 ;
        RECT 20.150 18.040 20.570 18.250 ;
        RECT 21.080 18.040 21.500 18.250 ;
        RECT 16.980 17.600 18.560 17.770 ;
        RECT 19.770 17.650 19.940 17.980 ;
        RECT 13.810 16.830 13.980 17.160 ;
        RECT 15.220 17.040 16.800 17.210 ;
        RECT 12.280 16.560 12.700 16.770 ;
        RECT 13.170 16.560 13.590 16.770 ;
        RECT 14.400 16.600 15.860 16.770 ;
        RECT 12.350 16.500 12.610 16.560 ;
        RECT 13.260 16.500 13.520 16.560 ;
        RECT 14.860 16.540 15.150 16.600 ;
        RECT 16.380 16.430 16.800 16.770 ;
        RECT 17.060 16.730 17.230 17.600 ;
        RECT 17.610 16.730 17.780 17.420 ;
        RECT 21.750 17.380 21.920 18.070 ;
        RECT 22.290 17.210 22.460 18.080 ;
        RECT 22.730 18.040 23.150 18.320 ;
        RECT 24.370 18.210 24.540 18.540 ;
        RECT 25.990 18.250 26.250 18.340 ;
        RECT 26.900 18.250 27.160 18.340 ;
        RECT 23.670 18.040 25.090 18.210 ;
        RECT 25.900 18.040 26.320 18.250 ;
        RECT 26.830 18.040 27.250 18.250 ;
        RECT 22.730 17.600 24.310 17.770 ;
        RECT 25.520 17.650 25.690 17.980 ;
        RECT 19.560 16.830 19.730 17.160 ;
        RECT 20.970 17.040 22.550 17.210 ;
        RECT 18.030 16.560 18.450 16.770 ;
        RECT 18.920 16.560 19.340 16.770 ;
        RECT 20.150 16.600 21.610 16.770 ;
        RECT 18.100 16.500 18.360 16.560 ;
        RECT 19.010 16.500 19.270 16.560 ;
        RECT 20.610 16.540 20.900 16.600 ;
        RECT 22.130 16.430 22.550 16.770 ;
        RECT 22.810 16.730 22.980 17.600 ;
        RECT 23.360 16.730 23.530 17.420 ;
        RECT 27.500 17.380 27.670 18.070 ;
        RECT 28.040 17.210 28.210 18.080 ;
        RECT 28.480 18.040 28.900 18.320 ;
        RECT 30.120 18.210 30.290 18.540 ;
        RECT 31.740 18.250 32.000 18.340 ;
        RECT 32.650 18.250 32.910 18.340 ;
        RECT 29.420 18.040 30.840 18.210 ;
        RECT 31.650 18.040 32.070 18.250 ;
        RECT 32.580 18.040 33.000 18.250 ;
        RECT 28.480 17.600 30.060 17.770 ;
        RECT 31.270 17.650 31.440 17.980 ;
        RECT 25.310 16.830 25.480 17.160 ;
        RECT 26.720 17.040 28.300 17.210 ;
        RECT 23.780 16.560 24.200 16.770 ;
        RECT 24.670 16.560 25.090 16.770 ;
        RECT 25.900 16.600 27.360 16.770 ;
        RECT 23.850 16.500 24.110 16.560 ;
        RECT 24.760 16.500 25.020 16.560 ;
        RECT 26.360 16.540 26.650 16.600 ;
        RECT 27.880 16.430 28.300 16.770 ;
        RECT 28.560 16.730 28.730 17.600 ;
        RECT 29.110 16.730 29.280 17.420 ;
        RECT 33.250 17.380 33.420 18.070 ;
        RECT 33.790 17.210 33.960 18.080 ;
        RECT 34.230 18.040 34.650 18.320 ;
        RECT 35.870 18.210 36.040 18.540 ;
        RECT 37.490 18.250 37.750 18.340 ;
        RECT 38.400 18.250 38.660 18.340 ;
        RECT 35.170 18.040 36.590 18.210 ;
        RECT 37.400 18.040 37.820 18.250 ;
        RECT 38.330 18.040 38.750 18.250 ;
        RECT 34.230 17.600 35.810 17.770 ;
        RECT 37.020 17.650 37.190 17.980 ;
        RECT 31.060 16.830 31.230 17.160 ;
        RECT 32.470 17.040 34.050 17.210 ;
        RECT 29.530 16.560 29.950 16.770 ;
        RECT 30.420 16.560 30.840 16.770 ;
        RECT 31.650 16.600 33.110 16.770 ;
        RECT 29.600 16.500 29.860 16.560 ;
        RECT 30.510 16.500 30.770 16.560 ;
        RECT 32.110 16.540 32.400 16.600 ;
        RECT 33.630 16.430 34.050 16.770 ;
        RECT 34.310 16.730 34.480 17.600 ;
        RECT 34.860 16.730 35.030 17.420 ;
        RECT 39.000 17.380 39.170 18.070 ;
        RECT 39.540 17.210 39.710 18.080 ;
        RECT 39.980 18.040 40.400 18.320 ;
        RECT 41.620 18.210 41.790 18.540 ;
        RECT 43.240 18.250 43.500 18.340 ;
        RECT 44.150 18.250 44.410 18.340 ;
        RECT 40.920 18.040 42.340 18.210 ;
        RECT 43.150 18.040 43.570 18.250 ;
        RECT 44.080 18.040 44.500 18.250 ;
        RECT 39.980 17.600 41.560 17.770 ;
        RECT 42.770 17.650 42.940 17.980 ;
        RECT 36.810 16.830 36.980 17.160 ;
        RECT 38.220 17.040 39.800 17.210 ;
        RECT 35.280 16.560 35.700 16.770 ;
        RECT 36.170 16.560 36.590 16.770 ;
        RECT 37.400 16.600 38.860 16.770 ;
        RECT 35.350 16.500 35.610 16.560 ;
        RECT 36.260 16.500 36.520 16.560 ;
        RECT 37.860 16.540 38.150 16.600 ;
        RECT 39.380 16.430 39.800 16.770 ;
        RECT 40.060 16.730 40.230 17.600 ;
        RECT 40.610 16.730 40.780 17.420 ;
        RECT 44.750 17.380 44.920 18.070 ;
        RECT 45.290 17.210 45.460 18.080 ;
        RECT 45.730 18.040 46.150 18.320 ;
        RECT 47.370 18.210 47.540 18.540 ;
        RECT 48.990 18.250 49.250 18.340 ;
        RECT 49.900 18.250 50.160 18.340 ;
        RECT 46.670 18.040 48.090 18.210 ;
        RECT 48.900 18.040 49.320 18.250 ;
        RECT 49.830 18.040 50.250 18.250 ;
        RECT 45.730 17.600 47.310 17.770 ;
        RECT 48.520 17.650 48.690 17.980 ;
        RECT 42.560 16.830 42.730 17.160 ;
        RECT 43.970 17.040 45.550 17.210 ;
        RECT 41.030 16.560 41.450 16.770 ;
        RECT 41.920 16.560 42.340 16.770 ;
        RECT 43.150 16.600 44.610 16.770 ;
        RECT 41.100 16.500 41.360 16.560 ;
        RECT 42.010 16.500 42.270 16.560 ;
        RECT 43.610 16.540 43.900 16.600 ;
        RECT 45.130 16.430 45.550 16.770 ;
        RECT 45.810 16.730 45.980 17.600 ;
        RECT 46.360 16.730 46.530 17.420 ;
        RECT 50.500 17.380 50.670 18.070 ;
        RECT 51.040 17.210 51.210 18.080 ;
        RECT 51.480 18.040 51.900 18.320 ;
        RECT 53.120 18.210 53.290 18.540 ;
        RECT 54.740 18.250 55.000 18.340 ;
        RECT 55.650 18.250 55.910 18.340 ;
        RECT 52.420 18.040 53.840 18.210 ;
        RECT 54.650 18.040 55.070 18.250 ;
        RECT 55.580 18.040 56.000 18.250 ;
        RECT 51.480 17.600 53.060 17.770 ;
        RECT 54.270 17.650 54.440 17.980 ;
        RECT 48.310 16.830 48.480 17.160 ;
        RECT 49.720 17.040 51.300 17.210 ;
        RECT 46.780 16.560 47.200 16.770 ;
        RECT 47.670 16.560 48.090 16.770 ;
        RECT 48.900 16.600 50.360 16.770 ;
        RECT 46.850 16.500 47.110 16.560 ;
        RECT 47.760 16.500 48.020 16.560 ;
        RECT 49.360 16.540 49.650 16.600 ;
        RECT 50.880 16.430 51.300 16.770 ;
        RECT 51.560 16.730 51.730 17.600 ;
        RECT 52.110 16.730 52.280 17.420 ;
        RECT 56.250 17.380 56.420 18.070 ;
        RECT 56.790 17.210 56.960 18.080 ;
        RECT 57.230 18.040 57.650 18.320 ;
        RECT 58.870 18.210 59.040 18.540 ;
        RECT 60.490 18.250 60.750 18.340 ;
        RECT 61.400 18.250 61.660 18.340 ;
        RECT 58.170 18.040 59.590 18.210 ;
        RECT 60.400 18.040 60.820 18.250 ;
        RECT 61.330 18.040 61.750 18.250 ;
        RECT 57.230 17.600 58.810 17.770 ;
        RECT 60.020 17.650 60.190 17.980 ;
        RECT 54.060 16.830 54.230 17.160 ;
        RECT 55.470 17.040 57.050 17.210 ;
        RECT 52.530 16.560 52.950 16.770 ;
        RECT 53.420 16.560 53.840 16.770 ;
        RECT 54.650 16.600 56.110 16.770 ;
        RECT 52.600 16.500 52.860 16.560 ;
        RECT 53.510 16.500 53.770 16.560 ;
        RECT 55.110 16.540 55.400 16.600 ;
        RECT 56.630 16.430 57.050 16.770 ;
        RECT 57.310 16.730 57.480 17.600 ;
        RECT 57.860 16.730 58.030 17.420 ;
        RECT 62.000 17.380 62.170 18.070 ;
        RECT 62.540 17.210 62.710 18.080 ;
        RECT 62.980 18.040 63.400 18.320 ;
        RECT 64.620 18.210 64.790 18.540 ;
        RECT 66.240 18.250 66.500 18.340 ;
        RECT 67.150 18.250 67.410 18.340 ;
        RECT 63.920 18.040 65.340 18.210 ;
        RECT 66.150 18.040 66.570 18.250 ;
        RECT 67.080 18.040 67.500 18.250 ;
        RECT 62.980 17.600 64.560 17.770 ;
        RECT 65.770 17.650 65.940 17.980 ;
        RECT 59.810 16.830 59.980 17.160 ;
        RECT 61.220 17.040 62.800 17.210 ;
        RECT 58.280 16.560 58.700 16.770 ;
        RECT 59.170 16.560 59.590 16.770 ;
        RECT 60.400 16.600 61.860 16.770 ;
        RECT 58.350 16.500 58.610 16.560 ;
        RECT 59.260 16.500 59.520 16.560 ;
        RECT 60.860 16.540 61.150 16.600 ;
        RECT 62.380 16.430 62.800 16.770 ;
        RECT 63.060 16.730 63.230 17.600 ;
        RECT 63.610 16.730 63.780 17.420 ;
        RECT 67.750 17.380 67.920 18.070 ;
        RECT 68.290 17.210 68.460 18.080 ;
        RECT 68.730 18.040 69.150 18.320 ;
        RECT 70.370 18.210 70.540 18.540 ;
        RECT 71.990 18.250 72.250 18.340 ;
        RECT 72.900 18.250 73.160 18.340 ;
        RECT 69.670 18.040 71.090 18.210 ;
        RECT 71.900 18.040 72.320 18.250 ;
        RECT 72.830 18.040 73.250 18.250 ;
        RECT 68.730 17.600 70.310 17.770 ;
        RECT 71.520 17.650 71.690 17.980 ;
        RECT 65.560 16.830 65.730 17.160 ;
        RECT 66.970 17.040 68.550 17.210 ;
        RECT 64.030 16.560 64.450 16.770 ;
        RECT 64.920 16.560 65.340 16.770 ;
        RECT 66.150 16.600 67.610 16.770 ;
        RECT 64.100 16.500 64.360 16.560 ;
        RECT 65.010 16.500 65.270 16.560 ;
        RECT 66.610 16.540 66.900 16.600 ;
        RECT 68.130 16.430 68.550 16.770 ;
        RECT 68.810 16.730 68.980 17.600 ;
        RECT 69.360 16.730 69.530 17.420 ;
        RECT 73.500 17.380 73.670 18.070 ;
        RECT 74.040 17.210 74.210 18.080 ;
        RECT 74.480 18.040 74.900 18.320 ;
        RECT 76.120 18.210 76.290 18.540 ;
        RECT 77.740 18.250 78.000 18.340 ;
        RECT 78.650 18.250 78.910 18.340 ;
        RECT 75.420 18.040 76.840 18.210 ;
        RECT 77.650 18.040 78.070 18.250 ;
        RECT 78.580 18.040 79.000 18.250 ;
        RECT 74.480 17.600 76.060 17.770 ;
        RECT 77.270 17.650 77.440 17.980 ;
        RECT 71.310 16.830 71.480 17.160 ;
        RECT 72.720 17.040 74.300 17.210 ;
        RECT 69.780 16.560 70.200 16.770 ;
        RECT 70.670 16.560 71.090 16.770 ;
        RECT 71.900 16.600 73.360 16.770 ;
        RECT 69.850 16.500 70.110 16.560 ;
        RECT 70.760 16.500 71.020 16.560 ;
        RECT 72.360 16.540 72.650 16.600 ;
        RECT 73.880 16.430 74.300 16.770 ;
        RECT 74.560 16.730 74.730 17.600 ;
        RECT 75.110 16.730 75.280 17.420 ;
        RECT 79.250 17.380 79.420 18.070 ;
        RECT 79.790 17.210 79.960 18.080 ;
        RECT 80.230 18.040 80.650 18.320 ;
        RECT 81.870 18.210 82.040 18.540 ;
        RECT 83.490 18.250 83.750 18.340 ;
        RECT 84.400 18.250 84.660 18.340 ;
        RECT 81.170 18.040 82.590 18.210 ;
        RECT 83.400 18.040 83.820 18.250 ;
        RECT 84.330 18.040 84.750 18.250 ;
        RECT 80.230 17.600 81.810 17.770 ;
        RECT 83.020 17.650 83.190 17.980 ;
        RECT 77.060 16.830 77.230 17.160 ;
        RECT 78.470 17.040 80.050 17.210 ;
        RECT 75.530 16.560 75.950 16.770 ;
        RECT 76.420 16.560 76.840 16.770 ;
        RECT 77.650 16.600 79.110 16.770 ;
        RECT 75.600 16.500 75.860 16.560 ;
        RECT 76.510 16.500 76.770 16.560 ;
        RECT 78.110 16.540 78.400 16.600 ;
        RECT 79.630 16.430 80.050 16.770 ;
        RECT 80.310 16.730 80.480 17.600 ;
        RECT 80.860 16.730 81.030 17.420 ;
        RECT 85.000 17.380 85.170 18.070 ;
        RECT 85.540 17.210 85.710 18.080 ;
        RECT 85.980 18.040 86.400 18.320 ;
        RECT 87.620 18.210 87.790 18.540 ;
        RECT 89.240 18.250 89.500 18.340 ;
        RECT 90.150 18.250 90.410 18.340 ;
        RECT 86.920 18.040 88.340 18.210 ;
        RECT 89.150 18.040 89.570 18.250 ;
        RECT 90.080 18.040 90.500 18.250 ;
        RECT 85.980 17.600 87.560 17.770 ;
        RECT 88.770 17.650 88.940 17.980 ;
        RECT 82.810 16.830 82.980 17.160 ;
        RECT 84.220 17.040 85.800 17.210 ;
        RECT 81.280 16.560 81.700 16.770 ;
        RECT 82.170 16.560 82.590 16.770 ;
        RECT 83.400 16.600 84.860 16.770 ;
        RECT 81.350 16.500 81.610 16.560 ;
        RECT 82.260 16.500 82.520 16.560 ;
        RECT 83.860 16.540 84.150 16.600 ;
        RECT 85.380 16.430 85.800 16.770 ;
        RECT 86.060 16.730 86.230 17.600 ;
        RECT 86.610 16.730 86.780 17.420 ;
        RECT 90.750 17.380 90.920 18.070 ;
        RECT 91.290 17.210 91.460 18.080 ;
        RECT 91.730 18.040 92.150 18.320 ;
        RECT 93.370 18.210 93.540 18.540 ;
        RECT 92.670 18.040 94.090 18.210 ;
        RECT 91.730 17.600 93.310 17.770 ;
        RECT 88.560 16.830 88.730 17.160 ;
        RECT 89.970 17.040 91.550 17.210 ;
        RECT 87.030 16.560 87.450 16.770 ;
        RECT 87.920 16.560 88.340 16.770 ;
        RECT 89.150 16.600 90.610 16.770 ;
        RECT 87.100 16.500 87.360 16.560 ;
        RECT 88.010 16.500 88.270 16.560 ;
        RECT 89.610 16.540 89.900 16.600 ;
        RECT 91.130 16.430 91.550 16.770 ;
        RECT 91.810 16.730 91.980 17.600 ;
        RECT 92.360 16.730 92.530 17.420 ;
        RECT 94.310 16.830 94.480 17.160 ;
        RECT 92.780 16.560 93.200 16.770 ;
        RECT 93.670 16.560 94.090 16.770 ;
        RECT 92.850 16.500 93.110 16.560 ;
        RECT 93.760 16.500 94.020 16.560 ;
        RECT 2.990 15.840 3.250 15.930 ;
        RECT 3.900 15.840 4.160 15.930 ;
        RECT 2.900 15.630 3.320 15.840 ;
        RECT 3.830 15.630 4.250 15.840 ;
        RECT 2.520 15.240 2.690 15.570 ;
        RECT 4.500 14.970 4.670 15.660 ;
        RECT 5.040 14.800 5.210 15.670 ;
        RECT 5.480 15.630 5.900 15.910 ;
        RECT 7.120 15.800 7.290 16.130 ;
        RECT 8.740 15.840 9.000 15.930 ;
        RECT 9.650 15.840 9.910 15.930 ;
        RECT 6.420 15.630 7.840 15.800 ;
        RECT 8.650 15.630 9.070 15.840 ;
        RECT 9.580 15.630 10.000 15.840 ;
        RECT 5.480 15.190 7.060 15.360 ;
        RECT 8.270 15.240 8.440 15.570 ;
        RECT 3.720 14.630 5.300 14.800 ;
        RECT 2.900 14.190 4.360 14.360 ;
        RECT 3.360 14.130 3.650 14.190 ;
        RECT 4.880 14.020 5.300 14.360 ;
        RECT 5.560 14.320 5.730 15.190 ;
        RECT 6.110 14.320 6.280 15.010 ;
        RECT 10.250 14.970 10.420 15.660 ;
        RECT 10.790 14.800 10.960 15.670 ;
        RECT 11.230 15.630 11.650 15.910 ;
        RECT 12.870 15.800 13.040 16.130 ;
        RECT 14.490 15.840 14.750 15.930 ;
        RECT 15.400 15.840 15.660 15.930 ;
        RECT 12.170 15.630 13.590 15.800 ;
        RECT 14.400 15.630 14.820 15.840 ;
        RECT 15.330 15.630 15.750 15.840 ;
        RECT 11.230 15.190 12.810 15.360 ;
        RECT 14.020 15.240 14.190 15.570 ;
        RECT 8.060 14.420 8.230 14.750 ;
        RECT 9.470 14.630 11.050 14.800 ;
        RECT 6.530 14.150 6.950 14.360 ;
        RECT 7.420 14.150 7.840 14.360 ;
        RECT 8.650 14.190 10.110 14.360 ;
        RECT 6.600 14.090 6.860 14.150 ;
        RECT 7.510 14.090 7.770 14.150 ;
        RECT 9.110 14.130 9.400 14.190 ;
        RECT 10.630 14.020 11.050 14.360 ;
        RECT 11.310 14.320 11.480 15.190 ;
        RECT 11.860 14.320 12.030 15.010 ;
        RECT 16.000 14.970 16.170 15.660 ;
        RECT 16.540 14.800 16.710 15.670 ;
        RECT 16.980 15.630 17.400 15.910 ;
        RECT 18.620 15.800 18.790 16.130 ;
        RECT 20.240 15.840 20.500 15.930 ;
        RECT 21.150 15.840 21.410 15.930 ;
        RECT 17.920 15.630 19.340 15.800 ;
        RECT 20.150 15.630 20.570 15.840 ;
        RECT 21.080 15.630 21.500 15.840 ;
        RECT 16.980 15.190 18.560 15.360 ;
        RECT 19.770 15.240 19.940 15.570 ;
        RECT 13.810 14.420 13.980 14.750 ;
        RECT 15.220 14.630 16.800 14.800 ;
        RECT 12.280 14.150 12.700 14.360 ;
        RECT 13.170 14.150 13.590 14.360 ;
        RECT 14.400 14.190 15.860 14.360 ;
        RECT 12.350 14.090 12.610 14.150 ;
        RECT 13.260 14.090 13.520 14.150 ;
        RECT 14.860 14.130 15.150 14.190 ;
        RECT 16.380 14.020 16.800 14.360 ;
        RECT 17.060 14.320 17.230 15.190 ;
        RECT 17.610 14.320 17.780 15.010 ;
        RECT 21.750 14.970 21.920 15.660 ;
        RECT 22.290 14.800 22.460 15.670 ;
        RECT 22.730 15.630 23.150 15.910 ;
        RECT 24.370 15.800 24.540 16.130 ;
        RECT 25.990 15.840 26.250 15.930 ;
        RECT 26.900 15.840 27.160 15.930 ;
        RECT 23.670 15.630 25.090 15.800 ;
        RECT 25.900 15.630 26.320 15.840 ;
        RECT 26.830 15.630 27.250 15.840 ;
        RECT 22.730 15.190 24.310 15.360 ;
        RECT 25.520 15.240 25.690 15.570 ;
        RECT 19.560 14.420 19.730 14.750 ;
        RECT 20.970 14.630 22.550 14.800 ;
        RECT 18.030 14.150 18.450 14.360 ;
        RECT 18.920 14.150 19.340 14.360 ;
        RECT 20.150 14.190 21.610 14.360 ;
        RECT 18.100 14.090 18.360 14.150 ;
        RECT 19.010 14.090 19.270 14.150 ;
        RECT 20.610 14.130 20.900 14.190 ;
        RECT 22.130 14.020 22.550 14.360 ;
        RECT 22.810 14.320 22.980 15.190 ;
        RECT 23.360 14.320 23.530 15.010 ;
        RECT 27.500 14.970 27.670 15.660 ;
        RECT 28.040 14.800 28.210 15.670 ;
        RECT 28.480 15.630 28.900 15.910 ;
        RECT 30.120 15.800 30.290 16.130 ;
        RECT 31.740 15.840 32.000 15.930 ;
        RECT 32.650 15.840 32.910 15.930 ;
        RECT 29.420 15.630 30.840 15.800 ;
        RECT 31.650 15.630 32.070 15.840 ;
        RECT 32.580 15.630 33.000 15.840 ;
        RECT 28.480 15.190 30.060 15.360 ;
        RECT 31.270 15.240 31.440 15.570 ;
        RECT 25.310 14.420 25.480 14.750 ;
        RECT 26.720 14.630 28.300 14.800 ;
        RECT 23.780 14.150 24.200 14.360 ;
        RECT 24.670 14.150 25.090 14.360 ;
        RECT 25.900 14.190 27.360 14.360 ;
        RECT 23.850 14.090 24.110 14.150 ;
        RECT 24.760 14.090 25.020 14.150 ;
        RECT 26.360 14.130 26.650 14.190 ;
        RECT 27.880 14.020 28.300 14.360 ;
        RECT 28.560 14.320 28.730 15.190 ;
        RECT 29.110 14.320 29.280 15.010 ;
        RECT 33.250 14.970 33.420 15.660 ;
        RECT 33.790 14.800 33.960 15.670 ;
        RECT 34.230 15.630 34.650 15.910 ;
        RECT 35.870 15.800 36.040 16.130 ;
        RECT 37.490 15.840 37.750 15.930 ;
        RECT 38.400 15.840 38.660 15.930 ;
        RECT 35.170 15.630 36.590 15.800 ;
        RECT 37.400 15.630 37.820 15.840 ;
        RECT 38.330 15.630 38.750 15.840 ;
        RECT 34.230 15.190 35.810 15.360 ;
        RECT 37.020 15.240 37.190 15.570 ;
        RECT 31.060 14.420 31.230 14.750 ;
        RECT 32.470 14.630 34.050 14.800 ;
        RECT 29.530 14.150 29.950 14.360 ;
        RECT 30.420 14.150 30.840 14.360 ;
        RECT 31.650 14.190 33.110 14.360 ;
        RECT 29.600 14.090 29.860 14.150 ;
        RECT 30.510 14.090 30.770 14.150 ;
        RECT 32.110 14.130 32.400 14.190 ;
        RECT 33.630 14.020 34.050 14.360 ;
        RECT 34.310 14.320 34.480 15.190 ;
        RECT 34.860 14.320 35.030 15.010 ;
        RECT 39.000 14.970 39.170 15.660 ;
        RECT 39.540 14.800 39.710 15.670 ;
        RECT 39.980 15.630 40.400 15.910 ;
        RECT 41.620 15.800 41.790 16.130 ;
        RECT 43.240 15.840 43.500 15.930 ;
        RECT 44.150 15.840 44.410 15.930 ;
        RECT 40.920 15.630 42.340 15.800 ;
        RECT 43.150 15.630 43.570 15.840 ;
        RECT 44.080 15.630 44.500 15.840 ;
        RECT 39.980 15.190 41.560 15.360 ;
        RECT 42.770 15.240 42.940 15.570 ;
        RECT 36.810 14.420 36.980 14.750 ;
        RECT 38.220 14.630 39.800 14.800 ;
        RECT 35.280 14.150 35.700 14.360 ;
        RECT 36.170 14.150 36.590 14.360 ;
        RECT 37.400 14.190 38.860 14.360 ;
        RECT 35.350 14.090 35.610 14.150 ;
        RECT 36.260 14.090 36.520 14.150 ;
        RECT 37.860 14.130 38.150 14.190 ;
        RECT 39.380 14.020 39.800 14.360 ;
        RECT 40.060 14.320 40.230 15.190 ;
        RECT 40.610 14.320 40.780 15.010 ;
        RECT 44.750 14.970 44.920 15.660 ;
        RECT 45.290 14.800 45.460 15.670 ;
        RECT 45.730 15.630 46.150 15.910 ;
        RECT 47.370 15.800 47.540 16.130 ;
        RECT 48.990 15.840 49.250 15.930 ;
        RECT 49.900 15.840 50.160 15.930 ;
        RECT 46.670 15.630 48.090 15.800 ;
        RECT 48.900 15.630 49.320 15.840 ;
        RECT 49.830 15.630 50.250 15.840 ;
        RECT 45.730 15.190 47.310 15.360 ;
        RECT 48.520 15.240 48.690 15.570 ;
        RECT 42.560 14.420 42.730 14.750 ;
        RECT 43.970 14.630 45.550 14.800 ;
        RECT 41.030 14.150 41.450 14.360 ;
        RECT 41.920 14.150 42.340 14.360 ;
        RECT 43.150 14.190 44.610 14.360 ;
        RECT 41.100 14.090 41.360 14.150 ;
        RECT 42.010 14.090 42.270 14.150 ;
        RECT 43.610 14.130 43.900 14.190 ;
        RECT 45.130 14.020 45.550 14.360 ;
        RECT 45.810 14.320 45.980 15.190 ;
        RECT 46.360 14.320 46.530 15.010 ;
        RECT 50.500 14.970 50.670 15.660 ;
        RECT 51.040 14.800 51.210 15.670 ;
        RECT 51.480 15.630 51.900 15.910 ;
        RECT 53.120 15.800 53.290 16.130 ;
        RECT 54.740 15.840 55.000 15.930 ;
        RECT 55.650 15.840 55.910 15.930 ;
        RECT 52.420 15.630 53.840 15.800 ;
        RECT 54.650 15.630 55.070 15.840 ;
        RECT 55.580 15.630 56.000 15.840 ;
        RECT 51.480 15.190 53.060 15.360 ;
        RECT 54.270 15.240 54.440 15.570 ;
        RECT 48.310 14.420 48.480 14.750 ;
        RECT 49.720 14.630 51.300 14.800 ;
        RECT 46.780 14.150 47.200 14.360 ;
        RECT 47.670 14.150 48.090 14.360 ;
        RECT 48.900 14.190 50.360 14.360 ;
        RECT 46.850 14.090 47.110 14.150 ;
        RECT 47.760 14.090 48.020 14.150 ;
        RECT 49.360 14.130 49.650 14.190 ;
        RECT 50.880 14.020 51.300 14.360 ;
        RECT 51.560 14.320 51.730 15.190 ;
        RECT 52.110 14.320 52.280 15.010 ;
        RECT 56.250 14.970 56.420 15.660 ;
        RECT 56.790 14.800 56.960 15.670 ;
        RECT 57.230 15.630 57.650 15.910 ;
        RECT 58.870 15.800 59.040 16.130 ;
        RECT 60.490 15.840 60.750 15.930 ;
        RECT 61.400 15.840 61.660 15.930 ;
        RECT 58.170 15.630 59.590 15.800 ;
        RECT 60.400 15.630 60.820 15.840 ;
        RECT 61.330 15.630 61.750 15.840 ;
        RECT 57.230 15.190 58.810 15.360 ;
        RECT 60.020 15.240 60.190 15.570 ;
        RECT 54.060 14.420 54.230 14.750 ;
        RECT 55.470 14.630 57.050 14.800 ;
        RECT 52.530 14.150 52.950 14.360 ;
        RECT 53.420 14.150 53.840 14.360 ;
        RECT 54.650 14.190 56.110 14.360 ;
        RECT 52.600 14.090 52.860 14.150 ;
        RECT 53.510 14.090 53.770 14.150 ;
        RECT 55.110 14.130 55.400 14.190 ;
        RECT 56.630 14.020 57.050 14.360 ;
        RECT 57.310 14.320 57.480 15.190 ;
        RECT 57.860 14.320 58.030 15.010 ;
        RECT 62.000 14.970 62.170 15.660 ;
        RECT 62.540 14.800 62.710 15.670 ;
        RECT 62.980 15.630 63.400 15.910 ;
        RECT 64.620 15.800 64.790 16.130 ;
        RECT 66.240 15.840 66.500 15.930 ;
        RECT 67.150 15.840 67.410 15.930 ;
        RECT 63.920 15.630 65.340 15.800 ;
        RECT 66.150 15.630 66.570 15.840 ;
        RECT 67.080 15.630 67.500 15.840 ;
        RECT 62.980 15.190 64.560 15.360 ;
        RECT 65.770 15.240 65.940 15.570 ;
        RECT 59.810 14.420 59.980 14.750 ;
        RECT 61.220 14.630 62.800 14.800 ;
        RECT 58.280 14.150 58.700 14.360 ;
        RECT 59.170 14.150 59.590 14.360 ;
        RECT 60.400 14.190 61.860 14.360 ;
        RECT 58.350 14.090 58.610 14.150 ;
        RECT 59.260 14.090 59.520 14.150 ;
        RECT 60.860 14.130 61.150 14.190 ;
        RECT 62.380 14.020 62.800 14.360 ;
        RECT 63.060 14.320 63.230 15.190 ;
        RECT 63.610 14.320 63.780 15.010 ;
        RECT 67.750 14.970 67.920 15.660 ;
        RECT 68.290 14.800 68.460 15.670 ;
        RECT 68.730 15.630 69.150 15.910 ;
        RECT 70.370 15.800 70.540 16.130 ;
        RECT 71.990 15.840 72.250 15.930 ;
        RECT 72.900 15.840 73.160 15.930 ;
        RECT 69.670 15.630 71.090 15.800 ;
        RECT 71.900 15.630 72.320 15.840 ;
        RECT 72.830 15.630 73.250 15.840 ;
        RECT 68.730 15.190 70.310 15.360 ;
        RECT 71.520 15.240 71.690 15.570 ;
        RECT 65.560 14.420 65.730 14.750 ;
        RECT 66.970 14.630 68.550 14.800 ;
        RECT 64.030 14.150 64.450 14.360 ;
        RECT 64.920 14.150 65.340 14.360 ;
        RECT 66.150 14.190 67.610 14.360 ;
        RECT 64.100 14.090 64.360 14.150 ;
        RECT 65.010 14.090 65.270 14.150 ;
        RECT 66.610 14.130 66.900 14.190 ;
        RECT 68.130 14.020 68.550 14.360 ;
        RECT 68.810 14.320 68.980 15.190 ;
        RECT 69.360 14.320 69.530 15.010 ;
        RECT 73.500 14.970 73.670 15.660 ;
        RECT 74.040 14.800 74.210 15.670 ;
        RECT 74.480 15.630 74.900 15.910 ;
        RECT 76.120 15.800 76.290 16.130 ;
        RECT 77.740 15.840 78.000 15.930 ;
        RECT 78.650 15.840 78.910 15.930 ;
        RECT 75.420 15.630 76.840 15.800 ;
        RECT 77.650 15.630 78.070 15.840 ;
        RECT 78.580 15.630 79.000 15.840 ;
        RECT 74.480 15.190 76.060 15.360 ;
        RECT 77.270 15.240 77.440 15.570 ;
        RECT 71.310 14.420 71.480 14.750 ;
        RECT 72.720 14.630 74.300 14.800 ;
        RECT 69.780 14.150 70.200 14.360 ;
        RECT 70.670 14.150 71.090 14.360 ;
        RECT 71.900 14.190 73.360 14.360 ;
        RECT 69.850 14.090 70.110 14.150 ;
        RECT 70.760 14.090 71.020 14.150 ;
        RECT 72.360 14.130 72.650 14.190 ;
        RECT 73.880 14.020 74.300 14.360 ;
        RECT 74.560 14.320 74.730 15.190 ;
        RECT 75.110 14.320 75.280 15.010 ;
        RECT 79.250 14.970 79.420 15.660 ;
        RECT 79.790 14.800 79.960 15.670 ;
        RECT 80.230 15.630 80.650 15.910 ;
        RECT 81.870 15.800 82.040 16.130 ;
        RECT 83.490 15.840 83.750 15.930 ;
        RECT 84.400 15.840 84.660 15.930 ;
        RECT 81.170 15.630 82.590 15.800 ;
        RECT 83.400 15.630 83.820 15.840 ;
        RECT 84.330 15.630 84.750 15.840 ;
        RECT 80.230 15.190 81.810 15.360 ;
        RECT 83.020 15.240 83.190 15.570 ;
        RECT 77.060 14.420 77.230 14.750 ;
        RECT 78.470 14.630 80.050 14.800 ;
        RECT 75.530 14.150 75.950 14.360 ;
        RECT 76.420 14.150 76.840 14.360 ;
        RECT 77.650 14.190 79.110 14.360 ;
        RECT 75.600 14.090 75.860 14.150 ;
        RECT 76.510 14.090 76.770 14.150 ;
        RECT 78.110 14.130 78.400 14.190 ;
        RECT 79.630 14.020 80.050 14.360 ;
        RECT 80.310 14.320 80.480 15.190 ;
        RECT 80.860 14.320 81.030 15.010 ;
        RECT 85.000 14.970 85.170 15.660 ;
        RECT 85.540 14.800 85.710 15.670 ;
        RECT 85.980 15.630 86.400 15.910 ;
        RECT 87.620 15.800 87.790 16.130 ;
        RECT 89.240 15.840 89.500 15.930 ;
        RECT 90.150 15.840 90.410 15.930 ;
        RECT 86.920 15.630 88.340 15.800 ;
        RECT 89.150 15.630 89.570 15.840 ;
        RECT 90.080 15.630 90.500 15.840 ;
        RECT 85.980 15.190 87.560 15.360 ;
        RECT 88.770 15.240 88.940 15.570 ;
        RECT 82.810 14.420 82.980 14.750 ;
        RECT 84.220 14.630 85.800 14.800 ;
        RECT 81.280 14.150 81.700 14.360 ;
        RECT 82.170 14.150 82.590 14.360 ;
        RECT 83.400 14.190 84.860 14.360 ;
        RECT 81.350 14.090 81.610 14.150 ;
        RECT 82.260 14.090 82.520 14.150 ;
        RECT 83.860 14.130 84.150 14.190 ;
        RECT 85.380 14.020 85.800 14.360 ;
        RECT 86.060 14.320 86.230 15.190 ;
        RECT 86.610 14.320 86.780 15.010 ;
        RECT 90.750 14.970 90.920 15.660 ;
        RECT 91.290 14.800 91.460 15.670 ;
        RECT 91.730 15.630 92.150 15.910 ;
        RECT 93.370 15.800 93.540 16.130 ;
        RECT 92.670 15.630 94.090 15.800 ;
        RECT 91.730 15.190 93.310 15.360 ;
        RECT 88.560 14.420 88.730 14.750 ;
        RECT 89.970 14.630 91.550 14.800 ;
        RECT 87.030 14.150 87.450 14.360 ;
        RECT 87.920 14.150 88.340 14.360 ;
        RECT 89.150 14.190 90.610 14.360 ;
        RECT 87.100 14.090 87.360 14.150 ;
        RECT 88.010 14.090 88.270 14.150 ;
        RECT 89.610 14.130 89.900 14.190 ;
        RECT 91.130 14.020 91.550 14.360 ;
        RECT 91.810 14.320 91.980 15.190 ;
        RECT 92.360 14.320 92.530 15.010 ;
        RECT 94.310 14.420 94.480 14.750 ;
        RECT 92.780 14.150 93.200 14.360 ;
        RECT 93.670 14.150 94.090 14.360 ;
        RECT 92.850 14.090 93.110 14.150 ;
        RECT 93.760 14.090 94.020 14.150 ;
        RECT 2.990 13.430 3.250 13.520 ;
        RECT 3.900 13.430 4.160 13.520 ;
        RECT 2.900 13.220 3.320 13.430 ;
        RECT 3.830 13.220 4.250 13.430 ;
        RECT 2.520 12.830 2.690 13.160 ;
        RECT 4.500 12.560 4.670 13.250 ;
        RECT 5.040 12.390 5.210 13.260 ;
        RECT 5.480 13.220 5.900 13.500 ;
        RECT 7.120 13.390 7.290 13.720 ;
        RECT 8.740 13.430 9.000 13.520 ;
        RECT 9.650 13.430 9.910 13.520 ;
        RECT 6.420 13.220 7.840 13.390 ;
        RECT 8.650 13.220 9.070 13.430 ;
        RECT 9.580 13.220 10.000 13.430 ;
        RECT 5.480 12.780 7.060 12.950 ;
        RECT 8.270 12.830 8.440 13.160 ;
        RECT 3.720 12.220 5.300 12.390 ;
        RECT 2.900 11.780 4.360 11.950 ;
        RECT 3.360 11.720 3.650 11.780 ;
        RECT 4.880 11.610 5.300 11.950 ;
        RECT 5.560 11.910 5.730 12.780 ;
        RECT 6.110 11.910 6.280 12.600 ;
        RECT 10.250 12.560 10.420 13.250 ;
        RECT 10.790 12.390 10.960 13.260 ;
        RECT 11.230 13.220 11.650 13.500 ;
        RECT 12.870 13.390 13.040 13.720 ;
        RECT 14.490 13.430 14.750 13.520 ;
        RECT 15.400 13.430 15.660 13.520 ;
        RECT 12.170 13.220 13.590 13.390 ;
        RECT 14.400 13.220 14.820 13.430 ;
        RECT 15.330 13.220 15.750 13.430 ;
        RECT 11.230 12.780 12.810 12.950 ;
        RECT 14.020 12.830 14.190 13.160 ;
        RECT 8.060 12.010 8.230 12.340 ;
        RECT 9.470 12.220 11.050 12.390 ;
        RECT 6.530 11.740 6.950 11.950 ;
        RECT 7.420 11.740 7.840 11.950 ;
        RECT 8.650 11.780 10.110 11.950 ;
        RECT 6.600 11.680 6.860 11.740 ;
        RECT 7.510 11.680 7.770 11.740 ;
        RECT 9.110 11.720 9.400 11.780 ;
        RECT 10.630 11.610 11.050 11.950 ;
        RECT 11.310 11.910 11.480 12.780 ;
        RECT 11.860 11.910 12.030 12.600 ;
        RECT 16.000 12.560 16.170 13.250 ;
        RECT 16.540 12.390 16.710 13.260 ;
        RECT 16.980 13.220 17.400 13.500 ;
        RECT 18.620 13.390 18.790 13.720 ;
        RECT 20.240 13.430 20.500 13.520 ;
        RECT 21.150 13.430 21.410 13.520 ;
        RECT 17.920 13.220 19.340 13.390 ;
        RECT 20.150 13.220 20.570 13.430 ;
        RECT 21.080 13.220 21.500 13.430 ;
        RECT 16.980 12.780 18.560 12.950 ;
        RECT 19.770 12.830 19.940 13.160 ;
        RECT 13.810 12.010 13.980 12.340 ;
        RECT 15.220 12.220 16.800 12.390 ;
        RECT 12.280 11.740 12.700 11.950 ;
        RECT 13.170 11.740 13.590 11.950 ;
        RECT 14.400 11.780 15.860 11.950 ;
        RECT 12.350 11.680 12.610 11.740 ;
        RECT 13.260 11.680 13.520 11.740 ;
        RECT 14.860 11.720 15.150 11.780 ;
        RECT 16.380 11.610 16.800 11.950 ;
        RECT 17.060 11.910 17.230 12.780 ;
        RECT 17.610 11.910 17.780 12.600 ;
        RECT 21.750 12.560 21.920 13.250 ;
        RECT 22.290 12.390 22.460 13.260 ;
        RECT 22.730 13.220 23.150 13.500 ;
        RECT 24.370 13.390 24.540 13.720 ;
        RECT 25.990 13.430 26.250 13.520 ;
        RECT 26.900 13.430 27.160 13.520 ;
        RECT 23.670 13.220 25.090 13.390 ;
        RECT 25.900 13.220 26.320 13.430 ;
        RECT 26.830 13.220 27.250 13.430 ;
        RECT 22.730 12.780 24.310 12.950 ;
        RECT 25.520 12.830 25.690 13.160 ;
        RECT 19.560 12.010 19.730 12.340 ;
        RECT 20.970 12.220 22.550 12.390 ;
        RECT 18.030 11.740 18.450 11.950 ;
        RECT 18.920 11.740 19.340 11.950 ;
        RECT 20.150 11.780 21.610 11.950 ;
        RECT 18.100 11.680 18.360 11.740 ;
        RECT 19.010 11.680 19.270 11.740 ;
        RECT 20.610 11.720 20.900 11.780 ;
        RECT 22.130 11.610 22.550 11.950 ;
        RECT 22.810 11.910 22.980 12.780 ;
        RECT 23.360 11.910 23.530 12.600 ;
        RECT 27.500 12.560 27.670 13.250 ;
        RECT 28.040 12.390 28.210 13.260 ;
        RECT 28.480 13.220 28.900 13.500 ;
        RECT 30.120 13.390 30.290 13.720 ;
        RECT 31.740 13.430 32.000 13.520 ;
        RECT 32.650 13.430 32.910 13.520 ;
        RECT 29.420 13.220 30.840 13.390 ;
        RECT 31.650 13.220 32.070 13.430 ;
        RECT 32.580 13.220 33.000 13.430 ;
        RECT 28.480 12.780 30.060 12.950 ;
        RECT 31.270 12.830 31.440 13.160 ;
        RECT 25.310 12.010 25.480 12.340 ;
        RECT 26.720 12.220 28.300 12.390 ;
        RECT 23.780 11.740 24.200 11.950 ;
        RECT 24.670 11.740 25.090 11.950 ;
        RECT 25.900 11.780 27.360 11.950 ;
        RECT 23.850 11.680 24.110 11.740 ;
        RECT 24.760 11.680 25.020 11.740 ;
        RECT 26.360 11.720 26.650 11.780 ;
        RECT 27.880 11.610 28.300 11.950 ;
        RECT 28.560 11.910 28.730 12.780 ;
        RECT 29.110 11.910 29.280 12.600 ;
        RECT 33.250 12.560 33.420 13.250 ;
        RECT 33.790 12.390 33.960 13.260 ;
        RECT 34.230 13.220 34.650 13.500 ;
        RECT 35.870 13.390 36.040 13.720 ;
        RECT 37.490 13.430 37.750 13.520 ;
        RECT 38.400 13.430 38.660 13.520 ;
        RECT 35.170 13.220 36.590 13.390 ;
        RECT 37.400 13.220 37.820 13.430 ;
        RECT 38.330 13.220 38.750 13.430 ;
        RECT 34.230 12.780 35.810 12.950 ;
        RECT 37.020 12.830 37.190 13.160 ;
        RECT 31.060 12.010 31.230 12.340 ;
        RECT 32.470 12.220 34.050 12.390 ;
        RECT 29.530 11.740 29.950 11.950 ;
        RECT 30.420 11.740 30.840 11.950 ;
        RECT 31.650 11.780 33.110 11.950 ;
        RECT 29.600 11.680 29.860 11.740 ;
        RECT 30.510 11.680 30.770 11.740 ;
        RECT 32.110 11.720 32.400 11.780 ;
        RECT 33.630 11.610 34.050 11.950 ;
        RECT 34.310 11.910 34.480 12.780 ;
        RECT 34.860 11.910 35.030 12.600 ;
        RECT 39.000 12.560 39.170 13.250 ;
        RECT 39.540 12.390 39.710 13.260 ;
        RECT 39.980 13.220 40.400 13.500 ;
        RECT 41.620 13.390 41.790 13.720 ;
        RECT 43.240 13.430 43.500 13.520 ;
        RECT 44.150 13.430 44.410 13.520 ;
        RECT 40.920 13.220 42.340 13.390 ;
        RECT 43.150 13.220 43.570 13.430 ;
        RECT 44.080 13.220 44.500 13.430 ;
        RECT 39.980 12.780 41.560 12.950 ;
        RECT 42.770 12.830 42.940 13.160 ;
        RECT 36.810 12.010 36.980 12.340 ;
        RECT 38.220 12.220 39.800 12.390 ;
        RECT 35.280 11.740 35.700 11.950 ;
        RECT 36.170 11.740 36.590 11.950 ;
        RECT 37.400 11.780 38.860 11.950 ;
        RECT 35.350 11.680 35.610 11.740 ;
        RECT 36.260 11.680 36.520 11.740 ;
        RECT 37.860 11.720 38.150 11.780 ;
        RECT 39.380 11.610 39.800 11.950 ;
        RECT 40.060 11.910 40.230 12.780 ;
        RECT 40.610 11.910 40.780 12.600 ;
        RECT 44.750 12.560 44.920 13.250 ;
        RECT 45.290 12.390 45.460 13.260 ;
        RECT 45.730 13.220 46.150 13.500 ;
        RECT 47.370 13.390 47.540 13.720 ;
        RECT 48.990 13.430 49.250 13.520 ;
        RECT 49.900 13.430 50.160 13.520 ;
        RECT 46.670 13.220 48.090 13.390 ;
        RECT 48.900 13.220 49.320 13.430 ;
        RECT 49.830 13.220 50.250 13.430 ;
        RECT 45.730 12.780 47.310 12.950 ;
        RECT 48.520 12.830 48.690 13.160 ;
        RECT 42.560 12.010 42.730 12.340 ;
        RECT 43.970 12.220 45.550 12.390 ;
        RECT 41.030 11.740 41.450 11.950 ;
        RECT 41.920 11.740 42.340 11.950 ;
        RECT 43.150 11.780 44.610 11.950 ;
        RECT 41.100 11.680 41.360 11.740 ;
        RECT 42.010 11.680 42.270 11.740 ;
        RECT 43.610 11.720 43.900 11.780 ;
        RECT 45.130 11.610 45.550 11.950 ;
        RECT 45.810 11.910 45.980 12.780 ;
        RECT 46.360 11.910 46.530 12.600 ;
        RECT 50.500 12.560 50.670 13.250 ;
        RECT 51.040 12.390 51.210 13.260 ;
        RECT 51.480 13.220 51.900 13.500 ;
        RECT 53.120 13.390 53.290 13.720 ;
        RECT 54.740 13.430 55.000 13.520 ;
        RECT 55.650 13.430 55.910 13.520 ;
        RECT 52.420 13.220 53.840 13.390 ;
        RECT 54.650 13.220 55.070 13.430 ;
        RECT 55.580 13.220 56.000 13.430 ;
        RECT 51.480 12.780 53.060 12.950 ;
        RECT 54.270 12.830 54.440 13.160 ;
        RECT 48.310 12.010 48.480 12.340 ;
        RECT 49.720 12.220 51.300 12.390 ;
        RECT 46.780 11.740 47.200 11.950 ;
        RECT 47.670 11.740 48.090 11.950 ;
        RECT 48.900 11.780 50.360 11.950 ;
        RECT 46.850 11.680 47.110 11.740 ;
        RECT 47.760 11.680 48.020 11.740 ;
        RECT 49.360 11.720 49.650 11.780 ;
        RECT 50.880 11.610 51.300 11.950 ;
        RECT 51.560 11.910 51.730 12.780 ;
        RECT 52.110 11.910 52.280 12.600 ;
        RECT 56.250 12.560 56.420 13.250 ;
        RECT 56.790 12.390 56.960 13.260 ;
        RECT 57.230 13.220 57.650 13.500 ;
        RECT 58.870 13.390 59.040 13.720 ;
        RECT 60.490 13.430 60.750 13.520 ;
        RECT 61.400 13.430 61.660 13.520 ;
        RECT 58.170 13.220 59.590 13.390 ;
        RECT 60.400 13.220 60.820 13.430 ;
        RECT 61.330 13.220 61.750 13.430 ;
        RECT 57.230 12.780 58.810 12.950 ;
        RECT 60.020 12.830 60.190 13.160 ;
        RECT 54.060 12.010 54.230 12.340 ;
        RECT 55.470 12.220 57.050 12.390 ;
        RECT 52.530 11.740 52.950 11.950 ;
        RECT 53.420 11.740 53.840 11.950 ;
        RECT 54.650 11.780 56.110 11.950 ;
        RECT 52.600 11.680 52.860 11.740 ;
        RECT 53.510 11.680 53.770 11.740 ;
        RECT 55.110 11.720 55.400 11.780 ;
        RECT 56.630 11.610 57.050 11.950 ;
        RECT 57.310 11.910 57.480 12.780 ;
        RECT 57.860 11.910 58.030 12.600 ;
        RECT 62.000 12.560 62.170 13.250 ;
        RECT 62.540 12.390 62.710 13.260 ;
        RECT 62.980 13.220 63.400 13.500 ;
        RECT 64.620 13.390 64.790 13.720 ;
        RECT 66.240 13.430 66.500 13.520 ;
        RECT 67.150 13.430 67.410 13.520 ;
        RECT 63.920 13.220 65.340 13.390 ;
        RECT 66.150 13.220 66.570 13.430 ;
        RECT 67.080 13.220 67.500 13.430 ;
        RECT 62.980 12.780 64.560 12.950 ;
        RECT 65.770 12.830 65.940 13.160 ;
        RECT 59.810 12.010 59.980 12.340 ;
        RECT 61.220 12.220 62.800 12.390 ;
        RECT 58.280 11.740 58.700 11.950 ;
        RECT 59.170 11.740 59.590 11.950 ;
        RECT 60.400 11.780 61.860 11.950 ;
        RECT 58.350 11.680 58.610 11.740 ;
        RECT 59.260 11.680 59.520 11.740 ;
        RECT 60.860 11.720 61.150 11.780 ;
        RECT 62.380 11.610 62.800 11.950 ;
        RECT 63.060 11.910 63.230 12.780 ;
        RECT 63.610 11.910 63.780 12.600 ;
        RECT 67.750 12.560 67.920 13.250 ;
        RECT 68.290 12.390 68.460 13.260 ;
        RECT 68.730 13.220 69.150 13.500 ;
        RECT 70.370 13.390 70.540 13.720 ;
        RECT 71.990 13.430 72.250 13.520 ;
        RECT 72.900 13.430 73.160 13.520 ;
        RECT 69.670 13.220 71.090 13.390 ;
        RECT 71.900 13.220 72.320 13.430 ;
        RECT 72.830 13.220 73.250 13.430 ;
        RECT 68.730 12.780 70.310 12.950 ;
        RECT 71.520 12.830 71.690 13.160 ;
        RECT 65.560 12.010 65.730 12.340 ;
        RECT 66.970 12.220 68.550 12.390 ;
        RECT 64.030 11.740 64.450 11.950 ;
        RECT 64.920 11.740 65.340 11.950 ;
        RECT 66.150 11.780 67.610 11.950 ;
        RECT 64.100 11.680 64.360 11.740 ;
        RECT 65.010 11.680 65.270 11.740 ;
        RECT 66.610 11.720 66.900 11.780 ;
        RECT 68.130 11.610 68.550 11.950 ;
        RECT 68.810 11.910 68.980 12.780 ;
        RECT 69.360 11.910 69.530 12.600 ;
        RECT 73.500 12.560 73.670 13.250 ;
        RECT 74.040 12.390 74.210 13.260 ;
        RECT 74.480 13.220 74.900 13.500 ;
        RECT 76.120 13.390 76.290 13.720 ;
        RECT 77.740 13.430 78.000 13.520 ;
        RECT 78.650 13.430 78.910 13.520 ;
        RECT 75.420 13.220 76.840 13.390 ;
        RECT 77.650 13.220 78.070 13.430 ;
        RECT 78.580 13.220 79.000 13.430 ;
        RECT 74.480 12.780 76.060 12.950 ;
        RECT 77.270 12.830 77.440 13.160 ;
        RECT 71.310 12.010 71.480 12.340 ;
        RECT 72.720 12.220 74.300 12.390 ;
        RECT 69.780 11.740 70.200 11.950 ;
        RECT 70.670 11.740 71.090 11.950 ;
        RECT 71.900 11.780 73.360 11.950 ;
        RECT 69.850 11.680 70.110 11.740 ;
        RECT 70.760 11.680 71.020 11.740 ;
        RECT 72.360 11.720 72.650 11.780 ;
        RECT 73.880 11.610 74.300 11.950 ;
        RECT 74.560 11.910 74.730 12.780 ;
        RECT 75.110 11.910 75.280 12.600 ;
        RECT 79.250 12.560 79.420 13.250 ;
        RECT 79.790 12.390 79.960 13.260 ;
        RECT 80.230 13.220 80.650 13.500 ;
        RECT 81.870 13.390 82.040 13.720 ;
        RECT 83.490 13.430 83.750 13.520 ;
        RECT 84.400 13.430 84.660 13.520 ;
        RECT 81.170 13.220 82.590 13.390 ;
        RECT 83.400 13.220 83.820 13.430 ;
        RECT 84.330 13.220 84.750 13.430 ;
        RECT 80.230 12.780 81.810 12.950 ;
        RECT 83.020 12.830 83.190 13.160 ;
        RECT 77.060 12.010 77.230 12.340 ;
        RECT 78.470 12.220 80.050 12.390 ;
        RECT 75.530 11.740 75.950 11.950 ;
        RECT 76.420 11.740 76.840 11.950 ;
        RECT 77.650 11.780 79.110 11.950 ;
        RECT 75.600 11.680 75.860 11.740 ;
        RECT 76.510 11.680 76.770 11.740 ;
        RECT 78.110 11.720 78.400 11.780 ;
        RECT 79.630 11.610 80.050 11.950 ;
        RECT 80.310 11.910 80.480 12.780 ;
        RECT 80.860 11.910 81.030 12.600 ;
        RECT 85.000 12.560 85.170 13.250 ;
        RECT 85.540 12.390 85.710 13.260 ;
        RECT 85.980 13.220 86.400 13.500 ;
        RECT 87.620 13.390 87.790 13.720 ;
        RECT 89.240 13.430 89.500 13.520 ;
        RECT 90.150 13.430 90.410 13.520 ;
        RECT 86.920 13.220 88.340 13.390 ;
        RECT 89.150 13.220 89.570 13.430 ;
        RECT 90.080 13.220 90.500 13.430 ;
        RECT 85.980 12.780 87.560 12.950 ;
        RECT 88.770 12.830 88.940 13.160 ;
        RECT 82.810 12.010 82.980 12.340 ;
        RECT 84.220 12.220 85.800 12.390 ;
        RECT 81.280 11.740 81.700 11.950 ;
        RECT 82.170 11.740 82.590 11.950 ;
        RECT 83.400 11.780 84.860 11.950 ;
        RECT 81.350 11.680 81.610 11.740 ;
        RECT 82.260 11.680 82.520 11.740 ;
        RECT 83.860 11.720 84.150 11.780 ;
        RECT 85.380 11.610 85.800 11.950 ;
        RECT 86.060 11.910 86.230 12.780 ;
        RECT 86.610 11.910 86.780 12.600 ;
        RECT 90.750 12.560 90.920 13.250 ;
        RECT 91.290 12.390 91.460 13.260 ;
        RECT 91.730 13.220 92.150 13.500 ;
        RECT 93.370 13.390 93.540 13.720 ;
        RECT 92.670 13.220 94.090 13.390 ;
        RECT 91.730 12.780 93.310 12.950 ;
        RECT 88.560 12.010 88.730 12.340 ;
        RECT 89.970 12.220 91.550 12.390 ;
        RECT 87.030 11.740 87.450 11.950 ;
        RECT 87.920 11.740 88.340 11.950 ;
        RECT 89.150 11.780 90.610 11.950 ;
        RECT 87.100 11.680 87.360 11.740 ;
        RECT 88.010 11.680 88.270 11.740 ;
        RECT 89.610 11.720 89.900 11.780 ;
        RECT 91.130 11.610 91.550 11.950 ;
        RECT 91.810 11.910 91.980 12.780 ;
        RECT 92.360 11.910 92.530 12.600 ;
        RECT 94.310 12.010 94.480 12.340 ;
        RECT 92.780 11.740 93.200 11.950 ;
        RECT 93.670 11.740 94.090 11.950 ;
        RECT 92.850 11.680 93.110 11.740 ;
        RECT 93.760 11.680 94.020 11.740 ;
        RECT 2.990 11.020 3.250 11.110 ;
        RECT 3.900 11.020 4.160 11.110 ;
        RECT 2.900 10.810 3.320 11.020 ;
        RECT 3.830 10.810 4.250 11.020 ;
        RECT 2.520 10.420 2.690 10.750 ;
        RECT 4.500 10.150 4.670 10.840 ;
        RECT 5.040 9.980 5.210 10.850 ;
        RECT 5.480 10.810 5.900 11.090 ;
        RECT 7.120 10.980 7.290 11.310 ;
        RECT 8.740 11.020 9.000 11.110 ;
        RECT 9.650 11.020 9.910 11.110 ;
        RECT 6.420 10.810 7.840 10.980 ;
        RECT 8.650 10.810 9.070 11.020 ;
        RECT 9.580 10.810 10.000 11.020 ;
        RECT 5.480 10.370 7.060 10.540 ;
        RECT 8.270 10.420 8.440 10.750 ;
        RECT 3.720 9.810 5.300 9.980 ;
        RECT 2.900 9.370 4.360 9.540 ;
        RECT 3.020 8.490 3.190 9.370 ;
        RECT 3.360 9.310 3.650 9.370 ;
        RECT 4.880 9.200 5.300 9.540 ;
        RECT 5.560 9.500 5.730 10.370 ;
        RECT 6.110 9.500 6.280 10.190 ;
        RECT 10.250 10.150 10.420 10.840 ;
        RECT 10.790 9.980 10.960 10.850 ;
        RECT 11.230 10.810 11.650 11.090 ;
        RECT 12.870 10.980 13.040 11.310 ;
        RECT 14.490 11.020 14.750 11.110 ;
        RECT 15.400 11.020 15.660 11.110 ;
        RECT 12.170 10.810 13.590 10.980 ;
        RECT 14.400 10.810 14.820 11.020 ;
        RECT 15.330 10.810 15.750 11.020 ;
        RECT 11.230 10.370 12.810 10.540 ;
        RECT 14.020 10.420 14.190 10.750 ;
        RECT 8.060 9.600 8.230 9.930 ;
        RECT 9.470 9.810 11.050 9.980 ;
        RECT 6.530 9.330 6.950 9.540 ;
        RECT 7.420 9.330 7.840 9.540 ;
        RECT 8.650 9.370 10.110 9.540 ;
        RECT 6.600 9.270 6.860 9.330 ;
        RECT 7.510 9.270 7.770 9.330 ;
        RECT 5.010 8.490 5.180 9.200 ;
        RECT 2.990 8.200 3.250 8.290 ;
        RECT 3.900 8.200 4.160 8.290 ;
        RECT 2.900 7.990 3.320 8.200 ;
        RECT 3.830 7.990 4.250 8.200 ;
        RECT 2.520 7.600 2.690 7.930 ;
        RECT 4.500 7.330 4.670 8.020 ;
        RECT 5.040 7.160 5.210 8.030 ;
        RECT 5.480 7.990 5.900 8.270 ;
        RECT 7.120 8.160 7.290 8.580 ;
        RECT 8.770 8.490 8.940 9.370 ;
        RECT 9.110 9.310 9.400 9.370 ;
        RECT 10.630 9.200 11.050 9.540 ;
        RECT 11.310 9.500 11.480 10.370 ;
        RECT 11.860 9.500 12.030 10.190 ;
        RECT 16.000 10.150 16.170 10.840 ;
        RECT 16.540 9.980 16.710 10.850 ;
        RECT 16.980 10.810 17.400 11.090 ;
        RECT 18.620 10.980 18.790 11.310 ;
        RECT 20.240 11.020 20.500 11.110 ;
        RECT 21.150 11.020 21.410 11.110 ;
        RECT 17.920 10.810 19.340 10.980 ;
        RECT 20.150 10.810 20.570 11.020 ;
        RECT 21.080 10.810 21.500 11.020 ;
        RECT 16.980 10.370 18.560 10.540 ;
        RECT 19.770 10.420 19.940 10.750 ;
        RECT 13.810 9.600 13.980 9.930 ;
        RECT 15.220 9.810 16.800 9.980 ;
        RECT 12.280 9.330 12.700 9.540 ;
        RECT 13.170 9.330 13.590 9.540 ;
        RECT 14.400 9.370 15.860 9.540 ;
        RECT 12.350 9.270 12.610 9.330 ;
        RECT 13.260 9.270 13.520 9.330 ;
        RECT 10.770 8.490 10.940 9.200 ;
        RECT 8.740 8.200 9.000 8.290 ;
        RECT 9.650 8.200 9.910 8.290 ;
        RECT 6.420 7.990 7.840 8.160 ;
        RECT 8.650 7.990 9.070 8.200 ;
        RECT 9.580 7.990 10.000 8.200 ;
        RECT 5.480 7.550 7.060 7.720 ;
        RECT 8.270 7.600 8.440 7.930 ;
        RECT 3.720 6.990 5.300 7.160 ;
        RECT 2.900 6.550 4.360 6.720 ;
        RECT 3.360 6.490 3.650 6.550 ;
        RECT 4.880 6.380 5.300 6.720 ;
        RECT 5.560 6.680 5.730 7.550 ;
        RECT 6.110 6.680 6.280 7.370 ;
        RECT 10.250 7.330 10.420 8.020 ;
        RECT 10.790 7.160 10.960 8.030 ;
        RECT 11.230 7.990 11.650 8.270 ;
        RECT 12.870 8.160 13.040 8.580 ;
        RECT 14.520 8.490 14.690 9.370 ;
        RECT 14.860 9.310 15.150 9.370 ;
        RECT 16.380 9.200 16.800 9.540 ;
        RECT 17.060 9.500 17.230 10.370 ;
        RECT 17.610 9.500 17.780 10.190 ;
        RECT 21.750 10.150 21.920 10.840 ;
        RECT 22.290 9.980 22.460 10.850 ;
        RECT 22.730 10.810 23.150 11.090 ;
        RECT 24.370 10.980 24.540 11.310 ;
        RECT 25.990 11.020 26.250 11.110 ;
        RECT 26.900 11.020 27.160 11.110 ;
        RECT 23.670 10.810 25.090 10.980 ;
        RECT 25.900 10.810 26.320 11.020 ;
        RECT 26.830 10.810 27.250 11.020 ;
        RECT 22.730 10.370 24.310 10.540 ;
        RECT 25.520 10.420 25.690 10.750 ;
        RECT 19.560 9.600 19.730 9.930 ;
        RECT 20.970 9.810 22.550 9.980 ;
        RECT 18.030 9.330 18.450 9.540 ;
        RECT 18.920 9.330 19.340 9.540 ;
        RECT 20.150 9.370 21.610 9.540 ;
        RECT 18.100 9.270 18.360 9.330 ;
        RECT 19.010 9.270 19.270 9.330 ;
        RECT 16.520 8.490 16.690 9.200 ;
        RECT 14.490 8.200 14.750 8.290 ;
        RECT 15.400 8.200 15.660 8.290 ;
        RECT 12.170 7.990 13.590 8.160 ;
        RECT 14.400 7.990 14.820 8.200 ;
        RECT 15.330 7.990 15.750 8.200 ;
        RECT 11.230 7.550 12.810 7.720 ;
        RECT 14.020 7.600 14.190 7.930 ;
        RECT 8.060 6.780 8.230 7.110 ;
        RECT 9.470 6.990 11.050 7.160 ;
        RECT 6.530 6.510 6.950 6.720 ;
        RECT 7.420 6.510 7.840 6.720 ;
        RECT 8.650 6.550 10.110 6.720 ;
        RECT 6.600 6.450 6.860 6.510 ;
        RECT 7.510 6.450 7.770 6.510 ;
        RECT 9.110 6.490 9.400 6.550 ;
        RECT 10.630 6.380 11.050 6.720 ;
        RECT 11.310 6.680 11.480 7.550 ;
        RECT 11.860 6.680 12.030 7.370 ;
        RECT 16.000 7.330 16.170 8.020 ;
        RECT 16.540 7.160 16.710 8.030 ;
        RECT 16.980 7.990 17.400 8.270 ;
        RECT 18.620 8.160 18.790 8.580 ;
        RECT 20.270 8.490 20.440 9.370 ;
        RECT 20.610 9.310 20.900 9.370 ;
        RECT 22.130 9.200 22.550 9.540 ;
        RECT 22.810 9.500 22.980 10.370 ;
        RECT 23.360 9.500 23.530 10.190 ;
        RECT 27.500 10.150 27.670 10.840 ;
        RECT 28.040 9.980 28.210 10.850 ;
        RECT 28.480 10.810 28.900 11.090 ;
        RECT 30.120 10.980 30.290 11.310 ;
        RECT 31.740 11.020 32.000 11.110 ;
        RECT 32.650 11.020 32.910 11.110 ;
        RECT 29.420 10.810 30.840 10.980 ;
        RECT 31.650 10.810 32.070 11.020 ;
        RECT 32.580 10.810 33.000 11.020 ;
        RECT 28.480 10.370 30.060 10.540 ;
        RECT 31.270 10.420 31.440 10.750 ;
        RECT 25.310 9.600 25.480 9.930 ;
        RECT 26.720 9.810 28.300 9.980 ;
        RECT 23.780 9.330 24.200 9.540 ;
        RECT 24.670 9.330 25.090 9.540 ;
        RECT 25.900 9.370 27.360 9.540 ;
        RECT 23.850 9.270 24.110 9.330 ;
        RECT 24.760 9.270 25.020 9.330 ;
        RECT 22.270 8.490 22.440 9.200 ;
        RECT 20.240 8.200 20.500 8.290 ;
        RECT 21.150 8.200 21.410 8.290 ;
        RECT 17.920 7.990 19.340 8.160 ;
        RECT 20.150 7.990 20.570 8.200 ;
        RECT 21.080 7.990 21.500 8.200 ;
        RECT 16.980 7.550 18.560 7.720 ;
        RECT 19.770 7.600 19.940 7.930 ;
        RECT 13.810 6.780 13.980 7.110 ;
        RECT 15.220 6.990 16.800 7.160 ;
        RECT 12.280 6.510 12.700 6.720 ;
        RECT 13.170 6.510 13.590 6.720 ;
        RECT 14.400 6.550 15.860 6.720 ;
        RECT 12.350 6.450 12.610 6.510 ;
        RECT 13.260 6.450 13.520 6.510 ;
        RECT 14.860 6.490 15.150 6.550 ;
        RECT 16.380 6.380 16.800 6.720 ;
        RECT 17.060 6.680 17.230 7.550 ;
        RECT 17.610 6.680 17.780 7.370 ;
        RECT 21.750 7.330 21.920 8.020 ;
        RECT 22.290 7.160 22.460 8.030 ;
        RECT 22.730 7.990 23.150 8.270 ;
        RECT 24.370 8.160 24.540 8.580 ;
        RECT 26.020 8.490 26.190 9.370 ;
        RECT 26.360 9.310 26.650 9.370 ;
        RECT 27.880 9.200 28.300 9.540 ;
        RECT 28.560 9.500 28.730 10.370 ;
        RECT 29.110 9.500 29.280 10.190 ;
        RECT 33.250 10.150 33.420 10.840 ;
        RECT 33.790 9.980 33.960 10.850 ;
        RECT 34.230 10.810 34.650 11.090 ;
        RECT 35.870 10.980 36.040 11.310 ;
        RECT 37.490 11.020 37.750 11.110 ;
        RECT 38.400 11.020 38.660 11.110 ;
        RECT 35.170 10.810 36.590 10.980 ;
        RECT 37.400 10.810 37.820 11.020 ;
        RECT 38.330 10.810 38.750 11.020 ;
        RECT 34.230 10.370 35.810 10.540 ;
        RECT 37.020 10.420 37.190 10.750 ;
        RECT 31.060 9.600 31.230 9.930 ;
        RECT 32.470 9.810 34.050 9.980 ;
        RECT 29.530 9.330 29.950 9.540 ;
        RECT 30.420 9.330 30.840 9.540 ;
        RECT 31.650 9.370 33.110 9.540 ;
        RECT 29.600 9.270 29.860 9.330 ;
        RECT 30.510 9.270 30.770 9.330 ;
        RECT 28.020 8.490 28.190 9.200 ;
        RECT 25.990 8.200 26.250 8.290 ;
        RECT 26.900 8.200 27.160 8.290 ;
        RECT 23.670 7.990 25.090 8.160 ;
        RECT 25.900 7.990 26.320 8.200 ;
        RECT 26.830 7.990 27.250 8.200 ;
        RECT 22.730 7.550 24.310 7.720 ;
        RECT 25.520 7.600 25.690 7.930 ;
        RECT 19.560 6.780 19.730 7.110 ;
        RECT 20.970 6.990 22.550 7.160 ;
        RECT 18.030 6.510 18.450 6.720 ;
        RECT 18.920 6.510 19.340 6.720 ;
        RECT 20.150 6.550 21.610 6.720 ;
        RECT 18.100 6.450 18.360 6.510 ;
        RECT 19.010 6.450 19.270 6.510 ;
        RECT 20.610 6.490 20.900 6.550 ;
        RECT 22.130 6.380 22.550 6.720 ;
        RECT 22.810 6.680 22.980 7.550 ;
        RECT 23.360 6.680 23.530 7.370 ;
        RECT 27.500 7.330 27.670 8.020 ;
        RECT 28.040 7.160 28.210 8.030 ;
        RECT 28.480 7.990 28.900 8.270 ;
        RECT 30.120 8.160 30.290 8.580 ;
        RECT 31.770 8.490 31.940 9.370 ;
        RECT 32.110 9.310 32.400 9.370 ;
        RECT 33.630 9.200 34.050 9.540 ;
        RECT 34.310 9.500 34.480 10.370 ;
        RECT 34.860 9.500 35.030 10.190 ;
        RECT 39.000 10.150 39.170 10.840 ;
        RECT 39.540 9.980 39.710 10.850 ;
        RECT 39.980 10.810 40.400 11.090 ;
        RECT 41.620 10.980 41.790 11.310 ;
        RECT 43.240 11.020 43.500 11.110 ;
        RECT 44.150 11.020 44.410 11.110 ;
        RECT 40.920 10.810 42.340 10.980 ;
        RECT 43.150 10.810 43.570 11.020 ;
        RECT 44.080 10.810 44.500 11.020 ;
        RECT 39.980 10.370 41.560 10.540 ;
        RECT 42.770 10.420 42.940 10.750 ;
        RECT 36.810 9.600 36.980 9.930 ;
        RECT 38.220 9.810 39.800 9.980 ;
        RECT 35.280 9.330 35.700 9.540 ;
        RECT 36.170 9.330 36.590 9.540 ;
        RECT 37.400 9.370 38.860 9.540 ;
        RECT 35.350 9.270 35.610 9.330 ;
        RECT 36.260 9.270 36.520 9.330 ;
        RECT 33.770 8.490 33.940 9.200 ;
        RECT 31.740 8.200 32.000 8.290 ;
        RECT 32.650 8.200 32.910 8.290 ;
        RECT 29.420 7.990 30.840 8.160 ;
        RECT 31.650 7.990 32.070 8.200 ;
        RECT 32.580 7.990 33.000 8.200 ;
        RECT 28.480 7.550 30.060 7.720 ;
        RECT 31.270 7.600 31.440 7.930 ;
        RECT 25.310 6.780 25.480 7.110 ;
        RECT 26.720 6.990 28.300 7.160 ;
        RECT 23.780 6.510 24.200 6.720 ;
        RECT 24.670 6.510 25.090 6.720 ;
        RECT 25.900 6.550 27.360 6.720 ;
        RECT 23.850 6.450 24.110 6.510 ;
        RECT 24.760 6.450 25.020 6.510 ;
        RECT 26.360 6.490 26.650 6.550 ;
        RECT 27.880 6.380 28.300 6.720 ;
        RECT 28.560 6.680 28.730 7.550 ;
        RECT 29.110 6.680 29.280 7.370 ;
        RECT 33.250 7.330 33.420 8.020 ;
        RECT 33.790 7.160 33.960 8.030 ;
        RECT 34.230 7.990 34.650 8.270 ;
        RECT 35.870 8.160 36.040 8.580 ;
        RECT 37.520 8.490 37.690 9.370 ;
        RECT 37.860 9.310 38.150 9.370 ;
        RECT 39.380 9.200 39.800 9.540 ;
        RECT 40.060 9.500 40.230 10.370 ;
        RECT 40.610 9.500 40.780 10.190 ;
        RECT 44.750 10.150 44.920 10.840 ;
        RECT 45.290 9.980 45.460 10.850 ;
        RECT 45.730 10.810 46.150 11.090 ;
        RECT 47.370 10.980 47.540 11.310 ;
        RECT 48.990 11.020 49.250 11.110 ;
        RECT 49.900 11.020 50.160 11.110 ;
        RECT 46.670 10.810 48.090 10.980 ;
        RECT 48.900 10.810 49.320 11.020 ;
        RECT 49.830 10.810 50.250 11.020 ;
        RECT 45.730 10.370 47.310 10.540 ;
        RECT 48.520 10.420 48.690 10.750 ;
        RECT 42.560 9.600 42.730 9.930 ;
        RECT 43.970 9.810 45.550 9.980 ;
        RECT 41.030 9.330 41.450 9.540 ;
        RECT 41.920 9.330 42.340 9.540 ;
        RECT 43.150 9.370 44.610 9.540 ;
        RECT 41.100 9.270 41.360 9.330 ;
        RECT 42.010 9.270 42.270 9.330 ;
        RECT 39.520 8.490 39.690 9.200 ;
        RECT 37.490 8.200 37.750 8.290 ;
        RECT 38.400 8.200 38.660 8.290 ;
        RECT 35.170 7.990 36.590 8.160 ;
        RECT 37.400 7.990 37.820 8.200 ;
        RECT 38.330 7.990 38.750 8.200 ;
        RECT 34.230 7.550 35.810 7.720 ;
        RECT 37.020 7.600 37.190 7.930 ;
        RECT 31.060 6.780 31.230 7.110 ;
        RECT 32.470 6.990 34.050 7.160 ;
        RECT 29.530 6.510 29.950 6.720 ;
        RECT 30.420 6.510 30.840 6.720 ;
        RECT 31.650 6.550 33.110 6.720 ;
        RECT 29.600 6.450 29.860 6.510 ;
        RECT 30.510 6.450 30.770 6.510 ;
        RECT 32.110 6.490 32.400 6.550 ;
        RECT 33.630 6.380 34.050 6.720 ;
        RECT 34.310 6.680 34.480 7.550 ;
        RECT 34.860 6.680 35.030 7.370 ;
        RECT 39.000 7.330 39.170 8.020 ;
        RECT 39.540 7.160 39.710 8.030 ;
        RECT 39.980 7.990 40.400 8.270 ;
        RECT 41.620 8.160 41.790 8.580 ;
        RECT 43.270 8.490 43.440 9.370 ;
        RECT 43.610 9.310 43.900 9.370 ;
        RECT 45.130 9.200 45.550 9.540 ;
        RECT 45.810 9.500 45.980 10.370 ;
        RECT 46.360 9.500 46.530 10.190 ;
        RECT 50.500 10.150 50.670 10.840 ;
        RECT 51.040 9.980 51.210 10.850 ;
        RECT 51.480 10.810 51.900 11.090 ;
        RECT 53.120 10.980 53.290 11.310 ;
        RECT 54.740 11.020 55.000 11.110 ;
        RECT 55.650 11.020 55.910 11.110 ;
        RECT 52.420 10.810 53.840 10.980 ;
        RECT 54.650 10.810 55.070 11.020 ;
        RECT 55.580 10.810 56.000 11.020 ;
        RECT 51.480 10.370 53.060 10.540 ;
        RECT 54.270 10.420 54.440 10.750 ;
        RECT 48.310 9.600 48.480 9.930 ;
        RECT 49.720 9.810 51.300 9.980 ;
        RECT 46.780 9.330 47.200 9.540 ;
        RECT 47.670 9.330 48.090 9.540 ;
        RECT 48.900 9.370 50.360 9.540 ;
        RECT 46.850 9.270 47.110 9.330 ;
        RECT 47.760 9.270 48.020 9.330 ;
        RECT 45.270 8.490 45.440 9.200 ;
        RECT 43.240 8.200 43.500 8.290 ;
        RECT 44.150 8.200 44.410 8.290 ;
        RECT 40.920 7.990 42.340 8.160 ;
        RECT 43.150 7.990 43.570 8.200 ;
        RECT 44.080 7.990 44.500 8.200 ;
        RECT 39.980 7.550 41.560 7.720 ;
        RECT 42.770 7.600 42.940 7.930 ;
        RECT 36.810 6.780 36.980 7.110 ;
        RECT 38.220 6.990 39.800 7.160 ;
        RECT 35.280 6.510 35.700 6.720 ;
        RECT 36.170 6.510 36.590 6.720 ;
        RECT 37.400 6.550 38.860 6.720 ;
        RECT 35.350 6.450 35.610 6.510 ;
        RECT 36.260 6.450 36.520 6.510 ;
        RECT 37.860 6.490 38.150 6.550 ;
        RECT 39.380 6.380 39.800 6.720 ;
        RECT 40.060 6.680 40.230 7.550 ;
        RECT 40.610 6.680 40.780 7.370 ;
        RECT 44.750 7.330 44.920 8.020 ;
        RECT 45.290 7.160 45.460 8.030 ;
        RECT 45.730 7.990 46.150 8.270 ;
        RECT 47.370 8.160 47.540 8.580 ;
        RECT 49.020 8.490 49.190 9.370 ;
        RECT 49.360 9.310 49.650 9.370 ;
        RECT 50.880 9.200 51.300 9.540 ;
        RECT 51.560 9.500 51.730 10.370 ;
        RECT 52.110 9.500 52.280 10.190 ;
        RECT 56.250 10.150 56.420 10.840 ;
        RECT 56.790 9.980 56.960 10.850 ;
        RECT 57.230 10.810 57.650 11.090 ;
        RECT 58.870 10.980 59.040 11.310 ;
        RECT 60.490 11.020 60.750 11.110 ;
        RECT 61.400 11.020 61.660 11.110 ;
        RECT 58.170 10.810 59.590 10.980 ;
        RECT 60.400 10.810 60.820 11.020 ;
        RECT 61.330 10.810 61.750 11.020 ;
        RECT 57.230 10.370 58.810 10.540 ;
        RECT 60.020 10.420 60.190 10.750 ;
        RECT 54.060 9.600 54.230 9.930 ;
        RECT 55.470 9.810 57.050 9.980 ;
        RECT 52.530 9.330 52.950 9.540 ;
        RECT 53.420 9.330 53.840 9.540 ;
        RECT 54.650 9.370 56.110 9.540 ;
        RECT 52.600 9.270 52.860 9.330 ;
        RECT 53.510 9.270 53.770 9.330 ;
        RECT 51.020 8.490 51.190 9.200 ;
        RECT 48.990 8.200 49.250 8.290 ;
        RECT 49.900 8.200 50.160 8.290 ;
        RECT 46.670 7.990 48.090 8.160 ;
        RECT 48.900 7.990 49.320 8.200 ;
        RECT 49.830 7.990 50.250 8.200 ;
        RECT 45.730 7.550 47.310 7.720 ;
        RECT 48.520 7.600 48.690 7.930 ;
        RECT 42.560 6.780 42.730 7.110 ;
        RECT 43.970 6.990 45.550 7.160 ;
        RECT 41.030 6.510 41.450 6.720 ;
        RECT 41.920 6.510 42.340 6.720 ;
        RECT 43.150 6.550 44.610 6.720 ;
        RECT 41.100 6.450 41.360 6.510 ;
        RECT 42.010 6.450 42.270 6.510 ;
        RECT 43.610 6.490 43.900 6.550 ;
        RECT 45.130 6.380 45.550 6.720 ;
        RECT 45.810 6.680 45.980 7.550 ;
        RECT 46.360 6.680 46.530 7.370 ;
        RECT 50.500 7.330 50.670 8.020 ;
        RECT 51.040 7.160 51.210 8.030 ;
        RECT 51.480 7.990 51.900 8.270 ;
        RECT 53.120 8.160 53.290 8.580 ;
        RECT 54.770 8.490 54.940 9.370 ;
        RECT 55.110 9.310 55.400 9.370 ;
        RECT 56.630 9.200 57.050 9.540 ;
        RECT 57.310 9.500 57.480 10.370 ;
        RECT 57.860 9.500 58.030 10.190 ;
        RECT 62.000 10.150 62.170 10.840 ;
        RECT 62.540 9.980 62.710 10.850 ;
        RECT 62.980 10.810 63.400 11.090 ;
        RECT 64.620 10.980 64.790 11.310 ;
        RECT 66.240 11.020 66.500 11.110 ;
        RECT 67.150 11.020 67.410 11.110 ;
        RECT 63.920 10.810 65.340 10.980 ;
        RECT 66.150 10.810 66.570 11.020 ;
        RECT 67.080 10.810 67.500 11.020 ;
        RECT 62.980 10.370 64.560 10.540 ;
        RECT 65.770 10.420 65.940 10.750 ;
        RECT 59.810 9.600 59.980 9.930 ;
        RECT 61.220 9.810 62.800 9.980 ;
        RECT 58.280 9.330 58.700 9.540 ;
        RECT 59.170 9.330 59.590 9.540 ;
        RECT 60.400 9.370 61.860 9.540 ;
        RECT 58.350 9.270 58.610 9.330 ;
        RECT 59.260 9.270 59.520 9.330 ;
        RECT 56.770 8.490 56.940 9.200 ;
        RECT 54.740 8.200 55.000 8.290 ;
        RECT 55.650 8.200 55.910 8.290 ;
        RECT 52.420 7.990 53.840 8.160 ;
        RECT 54.650 7.990 55.070 8.200 ;
        RECT 55.580 7.990 56.000 8.200 ;
        RECT 51.480 7.550 53.060 7.720 ;
        RECT 54.270 7.600 54.440 7.930 ;
        RECT 48.310 6.780 48.480 7.110 ;
        RECT 49.720 6.990 51.300 7.160 ;
        RECT 46.780 6.510 47.200 6.720 ;
        RECT 47.670 6.510 48.090 6.720 ;
        RECT 48.900 6.550 50.360 6.720 ;
        RECT 46.850 6.450 47.110 6.510 ;
        RECT 47.760 6.450 48.020 6.510 ;
        RECT 49.360 6.490 49.650 6.550 ;
        RECT 50.880 6.380 51.300 6.720 ;
        RECT 51.560 6.680 51.730 7.550 ;
        RECT 52.110 6.680 52.280 7.370 ;
        RECT 56.250 7.330 56.420 8.020 ;
        RECT 56.790 7.160 56.960 8.030 ;
        RECT 57.230 7.990 57.650 8.270 ;
        RECT 58.870 8.160 59.040 8.580 ;
        RECT 60.520 8.490 60.690 9.370 ;
        RECT 60.860 9.310 61.150 9.370 ;
        RECT 62.380 9.200 62.800 9.540 ;
        RECT 63.060 9.500 63.230 10.370 ;
        RECT 63.610 9.500 63.780 10.190 ;
        RECT 67.750 10.150 67.920 10.840 ;
        RECT 68.290 9.980 68.460 10.850 ;
        RECT 68.730 10.810 69.150 11.090 ;
        RECT 70.370 10.980 70.540 11.310 ;
        RECT 71.990 11.020 72.250 11.110 ;
        RECT 72.900 11.020 73.160 11.110 ;
        RECT 69.670 10.810 71.090 10.980 ;
        RECT 71.900 10.810 72.320 11.020 ;
        RECT 72.830 10.810 73.250 11.020 ;
        RECT 68.730 10.370 70.310 10.540 ;
        RECT 71.520 10.420 71.690 10.750 ;
        RECT 65.560 9.600 65.730 9.930 ;
        RECT 66.970 9.810 68.550 9.980 ;
        RECT 64.030 9.330 64.450 9.540 ;
        RECT 64.920 9.330 65.340 9.540 ;
        RECT 66.150 9.370 67.610 9.540 ;
        RECT 64.100 9.270 64.360 9.330 ;
        RECT 65.010 9.270 65.270 9.330 ;
        RECT 62.520 8.490 62.690 9.200 ;
        RECT 60.490 8.200 60.750 8.290 ;
        RECT 61.400 8.200 61.660 8.290 ;
        RECT 58.170 7.990 59.590 8.160 ;
        RECT 60.400 7.990 60.820 8.200 ;
        RECT 61.330 7.990 61.750 8.200 ;
        RECT 57.230 7.550 58.810 7.720 ;
        RECT 60.020 7.600 60.190 7.930 ;
        RECT 54.060 6.780 54.230 7.110 ;
        RECT 55.470 6.990 57.050 7.160 ;
        RECT 52.530 6.510 52.950 6.720 ;
        RECT 53.420 6.510 53.840 6.720 ;
        RECT 54.650 6.550 56.110 6.720 ;
        RECT 52.600 6.450 52.860 6.510 ;
        RECT 53.510 6.450 53.770 6.510 ;
        RECT 55.110 6.490 55.400 6.550 ;
        RECT 56.630 6.380 57.050 6.720 ;
        RECT 57.310 6.680 57.480 7.550 ;
        RECT 57.860 6.680 58.030 7.370 ;
        RECT 62.000 7.330 62.170 8.020 ;
        RECT 62.540 7.160 62.710 8.030 ;
        RECT 62.980 7.990 63.400 8.270 ;
        RECT 64.620 8.160 64.790 8.580 ;
        RECT 66.270 8.490 66.440 9.370 ;
        RECT 66.610 9.310 66.900 9.370 ;
        RECT 68.130 9.200 68.550 9.540 ;
        RECT 68.810 9.500 68.980 10.370 ;
        RECT 69.360 9.500 69.530 10.190 ;
        RECT 73.500 10.150 73.670 10.840 ;
        RECT 74.040 9.980 74.210 10.850 ;
        RECT 74.480 10.810 74.900 11.090 ;
        RECT 76.120 10.980 76.290 11.310 ;
        RECT 77.740 11.020 78.000 11.110 ;
        RECT 78.650 11.020 78.910 11.110 ;
        RECT 75.420 10.810 76.840 10.980 ;
        RECT 77.650 10.810 78.070 11.020 ;
        RECT 78.580 10.810 79.000 11.020 ;
        RECT 74.480 10.370 76.060 10.540 ;
        RECT 77.270 10.420 77.440 10.750 ;
        RECT 71.310 9.600 71.480 9.930 ;
        RECT 72.720 9.810 74.300 9.980 ;
        RECT 69.780 9.330 70.200 9.540 ;
        RECT 70.670 9.330 71.090 9.540 ;
        RECT 71.900 9.370 73.360 9.540 ;
        RECT 69.850 9.270 70.110 9.330 ;
        RECT 70.760 9.270 71.020 9.330 ;
        RECT 68.270 8.490 68.440 9.200 ;
        RECT 66.240 8.200 66.500 8.290 ;
        RECT 67.150 8.200 67.410 8.290 ;
        RECT 63.920 7.990 65.340 8.160 ;
        RECT 66.150 7.990 66.570 8.200 ;
        RECT 67.080 7.990 67.500 8.200 ;
        RECT 62.980 7.550 64.560 7.720 ;
        RECT 65.770 7.600 65.940 7.930 ;
        RECT 59.810 6.780 59.980 7.110 ;
        RECT 61.220 6.990 62.800 7.160 ;
        RECT 58.280 6.510 58.700 6.720 ;
        RECT 59.170 6.510 59.590 6.720 ;
        RECT 60.400 6.550 61.860 6.720 ;
        RECT 58.350 6.450 58.610 6.510 ;
        RECT 59.260 6.450 59.520 6.510 ;
        RECT 60.860 6.490 61.150 6.550 ;
        RECT 62.380 6.380 62.800 6.720 ;
        RECT 63.060 6.680 63.230 7.550 ;
        RECT 63.610 6.680 63.780 7.370 ;
        RECT 67.750 7.330 67.920 8.020 ;
        RECT 68.290 7.160 68.460 8.030 ;
        RECT 68.730 7.990 69.150 8.270 ;
        RECT 70.370 8.160 70.540 8.580 ;
        RECT 72.020 8.490 72.190 9.370 ;
        RECT 72.360 9.310 72.650 9.370 ;
        RECT 73.880 9.200 74.300 9.540 ;
        RECT 74.560 9.500 74.730 10.370 ;
        RECT 75.110 9.500 75.280 10.190 ;
        RECT 79.250 10.150 79.420 10.840 ;
        RECT 79.790 9.980 79.960 10.850 ;
        RECT 80.230 10.810 80.650 11.090 ;
        RECT 81.870 10.980 82.040 11.310 ;
        RECT 83.490 11.020 83.750 11.110 ;
        RECT 84.400 11.020 84.660 11.110 ;
        RECT 81.170 10.810 82.590 10.980 ;
        RECT 83.400 10.810 83.820 11.020 ;
        RECT 84.330 10.810 84.750 11.020 ;
        RECT 80.230 10.370 81.810 10.540 ;
        RECT 83.020 10.420 83.190 10.750 ;
        RECT 77.060 9.600 77.230 9.930 ;
        RECT 78.470 9.810 80.050 9.980 ;
        RECT 75.530 9.330 75.950 9.540 ;
        RECT 76.420 9.330 76.840 9.540 ;
        RECT 77.650 9.370 79.110 9.540 ;
        RECT 75.600 9.270 75.860 9.330 ;
        RECT 76.510 9.270 76.770 9.330 ;
        RECT 74.020 8.490 74.190 9.200 ;
        RECT 71.990 8.200 72.250 8.290 ;
        RECT 72.900 8.200 73.160 8.290 ;
        RECT 69.670 7.990 71.090 8.160 ;
        RECT 71.900 7.990 72.320 8.200 ;
        RECT 72.830 7.990 73.250 8.200 ;
        RECT 68.730 7.550 70.310 7.720 ;
        RECT 71.520 7.600 71.690 7.930 ;
        RECT 65.560 6.780 65.730 7.110 ;
        RECT 66.970 6.990 68.550 7.160 ;
        RECT 64.030 6.510 64.450 6.720 ;
        RECT 64.920 6.510 65.340 6.720 ;
        RECT 66.150 6.550 67.610 6.720 ;
        RECT 64.100 6.450 64.360 6.510 ;
        RECT 65.010 6.450 65.270 6.510 ;
        RECT 66.610 6.490 66.900 6.550 ;
        RECT 68.130 6.380 68.550 6.720 ;
        RECT 68.810 6.680 68.980 7.550 ;
        RECT 69.360 6.680 69.530 7.370 ;
        RECT 73.500 7.330 73.670 8.020 ;
        RECT 74.040 7.160 74.210 8.030 ;
        RECT 74.480 7.990 74.900 8.270 ;
        RECT 76.120 8.160 76.290 8.580 ;
        RECT 77.770 8.490 77.940 9.370 ;
        RECT 78.110 9.310 78.400 9.370 ;
        RECT 79.630 9.200 80.050 9.540 ;
        RECT 80.310 9.500 80.480 10.370 ;
        RECT 80.860 9.500 81.030 10.190 ;
        RECT 85.000 10.150 85.170 10.840 ;
        RECT 85.540 9.980 85.710 10.850 ;
        RECT 85.980 10.810 86.400 11.090 ;
        RECT 87.620 10.980 87.790 11.310 ;
        RECT 89.240 11.020 89.500 11.110 ;
        RECT 90.150 11.020 90.410 11.110 ;
        RECT 86.920 10.810 88.340 10.980 ;
        RECT 89.150 10.810 89.570 11.020 ;
        RECT 90.080 10.810 90.500 11.020 ;
        RECT 85.980 10.370 87.560 10.540 ;
        RECT 88.770 10.420 88.940 10.750 ;
        RECT 82.810 9.600 82.980 9.930 ;
        RECT 84.220 9.810 85.800 9.980 ;
        RECT 81.280 9.330 81.700 9.540 ;
        RECT 82.170 9.330 82.590 9.540 ;
        RECT 83.400 9.370 84.860 9.540 ;
        RECT 81.350 9.270 81.610 9.330 ;
        RECT 82.260 9.270 82.520 9.330 ;
        RECT 79.770 8.490 79.940 9.200 ;
        RECT 77.740 8.200 78.000 8.290 ;
        RECT 78.650 8.200 78.910 8.290 ;
        RECT 75.420 7.990 76.840 8.160 ;
        RECT 77.650 7.990 78.070 8.200 ;
        RECT 78.580 7.990 79.000 8.200 ;
        RECT 74.480 7.550 76.060 7.720 ;
        RECT 77.270 7.600 77.440 7.930 ;
        RECT 71.310 6.780 71.480 7.110 ;
        RECT 72.720 6.990 74.300 7.160 ;
        RECT 69.780 6.510 70.200 6.720 ;
        RECT 70.670 6.510 71.090 6.720 ;
        RECT 71.900 6.550 73.360 6.720 ;
        RECT 69.850 6.450 70.110 6.510 ;
        RECT 70.760 6.450 71.020 6.510 ;
        RECT 72.360 6.490 72.650 6.550 ;
        RECT 73.880 6.380 74.300 6.720 ;
        RECT 74.560 6.680 74.730 7.550 ;
        RECT 75.110 6.680 75.280 7.370 ;
        RECT 79.250 7.330 79.420 8.020 ;
        RECT 79.790 7.160 79.960 8.030 ;
        RECT 80.230 7.990 80.650 8.270 ;
        RECT 81.870 8.160 82.040 8.580 ;
        RECT 83.520 8.490 83.690 9.370 ;
        RECT 83.860 9.310 84.150 9.370 ;
        RECT 85.380 9.200 85.800 9.540 ;
        RECT 86.060 9.500 86.230 10.370 ;
        RECT 86.610 9.500 86.780 10.190 ;
        RECT 90.750 10.150 90.920 10.840 ;
        RECT 91.290 9.980 91.460 10.850 ;
        RECT 91.730 10.810 92.150 11.090 ;
        RECT 93.370 10.980 93.540 11.310 ;
        RECT 92.670 10.810 94.090 10.980 ;
        RECT 91.730 10.370 93.310 10.540 ;
        RECT 88.560 9.600 88.730 9.930 ;
        RECT 89.970 9.810 91.550 9.980 ;
        RECT 87.030 9.330 87.450 9.540 ;
        RECT 87.920 9.330 88.340 9.540 ;
        RECT 89.150 9.370 90.610 9.540 ;
        RECT 87.100 9.270 87.360 9.330 ;
        RECT 88.010 9.270 88.270 9.330 ;
        RECT 85.520 8.490 85.690 9.200 ;
        RECT 83.490 8.200 83.750 8.290 ;
        RECT 84.400 8.200 84.660 8.290 ;
        RECT 81.170 7.990 82.590 8.160 ;
        RECT 83.400 7.990 83.820 8.200 ;
        RECT 84.330 7.990 84.750 8.200 ;
        RECT 80.230 7.550 81.810 7.720 ;
        RECT 83.020 7.600 83.190 7.930 ;
        RECT 77.060 6.780 77.230 7.110 ;
        RECT 78.470 6.990 80.050 7.160 ;
        RECT 75.530 6.510 75.950 6.720 ;
        RECT 76.420 6.510 76.840 6.720 ;
        RECT 77.650 6.550 79.110 6.720 ;
        RECT 75.600 6.450 75.860 6.510 ;
        RECT 76.510 6.450 76.770 6.510 ;
        RECT 78.110 6.490 78.400 6.550 ;
        RECT 79.630 6.380 80.050 6.720 ;
        RECT 80.310 6.680 80.480 7.550 ;
        RECT 80.860 6.680 81.030 7.370 ;
        RECT 85.000 7.330 85.170 8.020 ;
        RECT 85.540 7.160 85.710 8.030 ;
        RECT 85.980 7.990 86.400 8.270 ;
        RECT 87.620 8.160 87.790 8.580 ;
        RECT 89.270 8.490 89.440 9.370 ;
        RECT 89.610 9.310 89.900 9.370 ;
        RECT 91.130 9.200 91.550 9.540 ;
        RECT 91.810 9.500 91.980 10.370 ;
        RECT 92.360 9.500 92.530 10.190 ;
        RECT 94.310 9.600 94.480 9.930 ;
        RECT 92.780 9.330 93.200 9.540 ;
        RECT 93.670 9.330 94.090 9.540 ;
        RECT 92.850 9.270 93.110 9.330 ;
        RECT 93.760 9.270 94.020 9.330 ;
        RECT 91.270 8.490 91.440 9.200 ;
        RECT 94.230 8.580 94.400 8.850 ;
        RECT 93.370 8.410 94.400 8.580 ;
        RECT 89.240 8.200 89.500 8.290 ;
        RECT 90.150 8.200 90.410 8.290 ;
        RECT 86.920 7.990 88.340 8.160 ;
        RECT 89.150 7.990 89.570 8.200 ;
        RECT 90.080 7.990 90.500 8.200 ;
        RECT 85.980 7.550 87.560 7.720 ;
        RECT 88.770 7.600 88.940 7.930 ;
        RECT 82.810 6.780 82.980 7.110 ;
        RECT 84.220 6.990 85.800 7.160 ;
        RECT 81.280 6.510 81.700 6.720 ;
        RECT 82.170 6.510 82.590 6.720 ;
        RECT 83.400 6.550 84.860 6.720 ;
        RECT 81.350 6.450 81.610 6.510 ;
        RECT 82.260 6.450 82.520 6.510 ;
        RECT 83.860 6.490 84.150 6.550 ;
        RECT 85.380 6.380 85.800 6.720 ;
        RECT 86.060 6.680 86.230 7.550 ;
        RECT 86.610 6.680 86.780 7.370 ;
        RECT 90.750 7.330 90.920 8.020 ;
        RECT 91.290 7.160 91.460 8.030 ;
        RECT 91.730 7.990 92.150 8.270 ;
        RECT 93.370 8.160 93.540 8.410 ;
        RECT 92.670 7.990 94.090 8.160 ;
        RECT 91.730 7.550 93.310 7.720 ;
        RECT 88.560 6.780 88.730 7.110 ;
        RECT 89.970 6.990 91.550 7.160 ;
        RECT 87.030 6.510 87.450 6.720 ;
        RECT 87.920 6.510 88.340 6.720 ;
        RECT 89.150 6.550 90.610 6.720 ;
        RECT 87.100 6.450 87.360 6.510 ;
        RECT 88.010 6.450 88.270 6.510 ;
        RECT 89.610 6.490 89.900 6.550 ;
        RECT 91.130 6.380 91.550 6.720 ;
        RECT 91.810 6.680 91.980 7.550 ;
        RECT 92.360 6.680 92.530 7.370 ;
        RECT 94.310 6.780 94.480 7.110 ;
        RECT 92.780 6.510 93.200 6.720 ;
        RECT 93.670 6.510 94.090 6.720 ;
        RECT 92.850 6.450 93.110 6.510 ;
        RECT 93.760 6.450 94.020 6.510 ;
        RECT 2.990 5.790 3.250 5.880 ;
        RECT 3.900 5.790 4.160 5.880 ;
        RECT 2.900 5.580 3.320 5.790 ;
        RECT 3.830 5.580 4.250 5.790 ;
        RECT 2.520 5.190 2.690 5.520 ;
        RECT 4.500 4.920 4.670 5.610 ;
        RECT 5.040 4.750 5.210 5.620 ;
        RECT 5.480 5.580 5.900 5.860 ;
        RECT 7.120 5.750 7.290 6.080 ;
        RECT 8.740 5.790 9.000 5.880 ;
        RECT 9.650 5.790 9.910 5.880 ;
        RECT 6.420 5.580 7.840 5.750 ;
        RECT 8.650 5.580 9.070 5.790 ;
        RECT 9.580 5.580 10.000 5.790 ;
        RECT 5.480 5.140 7.060 5.310 ;
        RECT 8.270 5.190 8.440 5.520 ;
        RECT 3.720 4.580 5.300 4.750 ;
        RECT 2.900 4.140 4.360 4.310 ;
        RECT 3.360 4.080 3.650 4.140 ;
        RECT 4.880 3.970 5.300 4.310 ;
        RECT 5.560 4.270 5.730 5.140 ;
        RECT 6.110 4.270 6.280 4.960 ;
        RECT 10.250 4.920 10.420 5.610 ;
        RECT 10.790 4.750 10.960 5.620 ;
        RECT 11.230 5.580 11.650 5.860 ;
        RECT 12.870 5.750 13.040 6.080 ;
        RECT 14.490 5.790 14.750 5.880 ;
        RECT 15.400 5.790 15.660 5.880 ;
        RECT 12.170 5.580 13.590 5.750 ;
        RECT 14.400 5.580 14.820 5.790 ;
        RECT 15.330 5.580 15.750 5.790 ;
        RECT 11.230 5.140 12.810 5.310 ;
        RECT 14.020 5.190 14.190 5.520 ;
        RECT 8.060 4.370 8.230 4.700 ;
        RECT 9.470 4.580 11.050 4.750 ;
        RECT 6.530 4.100 6.950 4.310 ;
        RECT 7.420 4.100 7.840 4.310 ;
        RECT 8.650 4.140 10.110 4.310 ;
        RECT 6.600 4.040 6.860 4.100 ;
        RECT 7.510 4.040 7.770 4.100 ;
        RECT 9.110 4.080 9.400 4.140 ;
        RECT 10.630 3.970 11.050 4.310 ;
        RECT 11.310 4.270 11.480 5.140 ;
        RECT 11.860 4.270 12.030 4.960 ;
        RECT 16.000 4.920 16.170 5.610 ;
        RECT 16.540 4.750 16.710 5.620 ;
        RECT 16.980 5.580 17.400 5.860 ;
        RECT 18.620 5.750 18.790 6.080 ;
        RECT 20.240 5.790 20.500 5.880 ;
        RECT 21.150 5.790 21.410 5.880 ;
        RECT 17.920 5.580 19.340 5.750 ;
        RECT 20.150 5.580 20.570 5.790 ;
        RECT 21.080 5.580 21.500 5.790 ;
        RECT 16.980 5.140 18.560 5.310 ;
        RECT 19.770 5.190 19.940 5.520 ;
        RECT 13.810 4.370 13.980 4.700 ;
        RECT 15.220 4.580 16.800 4.750 ;
        RECT 12.280 4.100 12.700 4.310 ;
        RECT 13.170 4.100 13.590 4.310 ;
        RECT 14.400 4.140 15.860 4.310 ;
        RECT 12.350 4.040 12.610 4.100 ;
        RECT 13.260 4.040 13.520 4.100 ;
        RECT 14.860 4.080 15.150 4.140 ;
        RECT 16.380 3.970 16.800 4.310 ;
        RECT 17.060 4.270 17.230 5.140 ;
        RECT 17.610 4.270 17.780 4.960 ;
        RECT 21.750 4.920 21.920 5.610 ;
        RECT 22.290 4.750 22.460 5.620 ;
        RECT 22.730 5.580 23.150 5.860 ;
        RECT 24.370 5.750 24.540 6.080 ;
        RECT 25.990 5.790 26.250 5.880 ;
        RECT 26.900 5.790 27.160 5.880 ;
        RECT 23.670 5.580 25.090 5.750 ;
        RECT 25.900 5.580 26.320 5.790 ;
        RECT 26.830 5.580 27.250 5.790 ;
        RECT 22.730 5.140 24.310 5.310 ;
        RECT 25.520 5.190 25.690 5.520 ;
        RECT 19.560 4.370 19.730 4.700 ;
        RECT 20.970 4.580 22.550 4.750 ;
        RECT 18.030 4.100 18.450 4.310 ;
        RECT 18.920 4.100 19.340 4.310 ;
        RECT 20.150 4.140 21.610 4.310 ;
        RECT 18.100 4.040 18.360 4.100 ;
        RECT 19.010 4.040 19.270 4.100 ;
        RECT 20.610 4.080 20.900 4.140 ;
        RECT 22.130 3.970 22.550 4.310 ;
        RECT 22.810 4.270 22.980 5.140 ;
        RECT 23.360 4.270 23.530 4.960 ;
        RECT 27.500 4.920 27.670 5.610 ;
        RECT 28.040 4.750 28.210 5.620 ;
        RECT 28.480 5.580 28.900 5.860 ;
        RECT 30.120 5.750 30.290 6.080 ;
        RECT 31.740 5.790 32.000 5.880 ;
        RECT 32.650 5.790 32.910 5.880 ;
        RECT 29.420 5.580 30.840 5.750 ;
        RECT 31.650 5.580 32.070 5.790 ;
        RECT 32.580 5.580 33.000 5.790 ;
        RECT 28.480 5.140 30.060 5.310 ;
        RECT 31.270 5.190 31.440 5.520 ;
        RECT 25.310 4.370 25.480 4.700 ;
        RECT 26.720 4.580 28.300 4.750 ;
        RECT 23.780 4.100 24.200 4.310 ;
        RECT 24.670 4.100 25.090 4.310 ;
        RECT 25.900 4.140 27.360 4.310 ;
        RECT 23.850 4.040 24.110 4.100 ;
        RECT 24.760 4.040 25.020 4.100 ;
        RECT 26.360 4.080 26.650 4.140 ;
        RECT 27.880 3.970 28.300 4.310 ;
        RECT 28.560 4.270 28.730 5.140 ;
        RECT 29.110 4.270 29.280 4.960 ;
        RECT 33.250 4.920 33.420 5.610 ;
        RECT 33.790 4.750 33.960 5.620 ;
        RECT 34.230 5.580 34.650 5.860 ;
        RECT 35.870 5.750 36.040 6.080 ;
        RECT 37.490 5.790 37.750 5.880 ;
        RECT 38.400 5.790 38.660 5.880 ;
        RECT 35.170 5.580 36.590 5.750 ;
        RECT 37.400 5.580 37.820 5.790 ;
        RECT 38.330 5.580 38.750 5.790 ;
        RECT 34.230 5.140 35.810 5.310 ;
        RECT 37.020 5.190 37.190 5.520 ;
        RECT 31.060 4.370 31.230 4.700 ;
        RECT 32.470 4.580 34.050 4.750 ;
        RECT 29.530 4.100 29.950 4.310 ;
        RECT 30.420 4.100 30.840 4.310 ;
        RECT 31.650 4.140 33.110 4.310 ;
        RECT 29.600 4.040 29.860 4.100 ;
        RECT 30.510 4.040 30.770 4.100 ;
        RECT 32.110 4.080 32.400 4.140 ;
        RECT 33.630 3.970 34.050 4.310 ;
        RECT 34.310 4.270 34.480 5.140 ;
        RECT 34.860 4.270 35.030 4.960 ;
        RECT 39.000 4.920 39.170 5.610 ;
        RECT 39.540 4.750 39.710 5.620 ;
        RECT 39.980 5.580 40.400 5.860 ;
        RECT 41.620 5.750 41.790 6.080 ;
        RECT 43.240 5.790 43.500 5.880 ;
        RECT 44.150 5.790 44.410 5.880 ;
        RECT 40.920 5.580 42.340 5.750 ;
        RECT 43.150 5.580 43.570 5.790 ;
        RECT 44.080 5.580 44.500 5.790 ;
        RECT 39.980 5.140 41.560 5.310 ;
        RECT 42.770 5.190 42.940 5.520 ;
        RECT 36.810 4.370 36.980 4.700 ;
        RECT 38.220 4.580 39.800 4.750 ;
        RECT 35.280 4.100 35.700 4.310 ;
        RECT 36.170 4.100 36.590 4.310 ;
        RECT 37.400 4.140 38.860 4.310 ;
        RECT 35.350 4.040 35.610 4.100 ;
        RECT 36.260 4.040 36.520 4.100 ;
        RECT 37.860 4.080 38.150 4.140 ;
        RECT 39.380 3.970 39.800 4.310 ;
        RECT 40.060 4.270 40.230 5.140 ;
        RECT 40.610 4.270 40.780 4.960 ;
        RECT 44.750 4.920 44.920 5.610 ;
        RECT 45.290 4.750 45.460 5.620 ;
        RECT 45.730 5.580 46.150 5.860 ;
        RECT 47.370 5.750 47.540 6.080 ;
        RECT 48.990 5.790 49.250 5.880 ;
        RECT 49.900 5.790 50.160 5.880 ;
        RECT 46.670 5.580 48.090 5.750 ;
        RECT 48.900 5.580 49.320 5.790 ;
        RECT 49.830 5.580 50.250 5.790 ;
        RECT 45.730 5.140 47.310 5.310 ;
        RECT 48.520 5.190 48.690 5.520 ;
        RECT 42.560 4.370 42.730 4.700 ;
        RECT 43.970 4.580 45.550 4.750 ;
        RECT 41.030 4.100 41.450 4.310 ;
        RECT 41.920 4.100 42.340 4.310 ;
        RECT 43.150 4.140 44.610 4.310 ;
        RECT 41.100 4.040 41.360 4.100 ;
        RECT 42.010 4.040 42.270 4.100 ;
        RECT 43.610 4.080 43.900 4.140 ;
        RECT 45.130 3.970 45.550 4.310 ;
        RECT 45.810 4.270 45.980 5.140 ;
        RECT 46.360 4.270 46.530 4.960 ;
        RECT 50.500 4.920 50.670 5.610 ;
        RECT 51.040 4.750 51.210 5.620 ;
        RECT 51.480 5.580 51.900 5.860 ;
        RECT 53.120 5.750 53.290 6.080 ;
        RECT 54.740 5.790 55.000 5.880 ;
        RECT 55.650 5.790 55.910 5.880 ;
        RECT 52.420 5.580 53.840 5.750 ;
        RECT 54.650 5.580 55.070 5.790 ;
        RECT 55.580 5.580 56.000 5.790 ;
        RECT 51.480 5.140 53.060 5.310 ;
        RECT 54.270 5.190 54.440 5.520 ;
        RECT 48.310 4.370 48.480 4.700 ;
        RECT 49.720 4.580 51.300 4.750 ;
        RECT 46.780 4.100 47.200 4.310 ;
        RECT 47.670 4.100 48.090 4.310 ;
        RECT 48.900 4.140 50.360 4.310 ;
        RECT 46.850 4.040 47.110 4.100 ;
        RECT 47.760 4.040 48.020 4.100 ;
        RECT 49.360 4.080 49.650 4.140 ;
        RECT 50.880 3.970 51.300 4.310 ;
        RECT 51.560 4.270 51.730 5.140 ;
        RECT 52.110 4.270 52.280 4.960 ;
        RECT 56.250 4.920 56.420 5.610 ;
        RECT 56.790 4.750 56.960 5.620 ;
        RECT 57.230 5.580 57.650 5.860 ;
        RECT 58.870 5.750 59.040 6.080 ;
        RECT 60.490 5.790 60.750 5.880 ;
        RECT 61.400 5.790 61.660 5.880 ;
        RECT 58.170 5.580 59.590 5.750 ;
        RECT 60.400 5.580 60.820 5.790 ;
        RECT 61.330 5.580 61.750 5.790 ;
        RECT 57.230 5.140 58.810 5.310 ;
        RECT 60.020 5.190 60.190 5.520 ;
        RECT 54.060 4.370 54.230 4.700 ;
        RECT 55.470 4.580 57.050 4.750 ;
        RECT 52.530 4.100 52.950 4.310 ;
        RECT 53.420 4.100 53.840 4.310 ;
        RECT 54.650 4.140 56.110 4.310 ;
        RECT 52.600 4.040 52.860 4.100 ;
        RECT 53.510 4.040 53.770 4.100 ;
        RECT 55.110 4.080 55.400 4.140 ;
        RECT 56.630 3.970 57.050 4.310 ;
        RECT 57.310 4.270 57.480 5.140 ;
        RECT 57.860 4.270 58.030 4.960 ;
        RECT 62.000 4.920 62.170 5.610 ;
        RECT 62.540 4.750 62.710 5.620 ;
        RECT 62.980 5.580 63.400 5.860 ;
        RECT 64.620 5.750 64.790 6.080 ;
        RECT 66.240 5.790 66.500 5.880 ;
        RECT 67.150 5.790 67.410 5.880 ;
        RECT 63.920 5.580 65.340 5.750 ;
        RECT 66.150 5.580 66.570 5.790 ;
        RECT 67.080 5.580 67.500 5.790 ;
        RECT 62.980 5.140 64.560 5.310 ;
        RECT 65.770 5.190 65.940 5.520 ;
        RECT 59.810 4.370 59.980 4.700 ;
        RECT 61.220 4.580 62.800 4.750 ;
        RECT 58.280 4.100 58.700 4.310 ;
        RECT 59.170 4.100 59.590 4.310 ;
        RECT 60.400 4.140 61.860 4.310 ;
        RECT 58.350 4.040 58.610 4.100 ;
        RECT 59.260 4.040 59.520 4.100 ;
        RECT 60.860 4.080 61.150 4.140 ;
        RECT 62.380 3.970 62.800 4.310 ;
        RECT 63.060 4.270 63.230 5.140 ;
        RECT 63.610 4.270 63.780 4.960 ;
        RECT 67.750 4.920 67.920 5.610 ;
        RECT 68.290 4.750 68.460 5.620 ;
        RECT 68.730 5.580 69.150 5.860 ;
        RECT 70.370 5.750 70.540 6.080 ;
        RECT 71.990 5.790 72.250 5.880 ;
        RECT 72.900 5.790 73.160 5.880 ;
        RECT 69.670 5.580 71.090 5.750 ;
        RECT 71.900 5.580 72.320 5.790 ;
        RECT 72.830 5.580 73.250 5.790 ;
        RECT 68.730 5.140 70.310 5.310 ;
        RECT 71.520 5.190 71.690 5.520 ;
        RECT 65.560 4.370 65.730 4.700 ;
        RECT 66.970 4.580 68.550 4.750 ;
        RECT 64.030 4.100 64.450 4.310 ;
        RECT 64.920 4.100 65.340 4.310 ;
        RECT 66.150 4.140 67.610 4.310 ;
        RECT 64.100 4.040 64.360 4.100 ;
        RECT 65.010 4.040 65.270 4.100 ;
        RECT 66.610 4.080 66.900 4.140 ;
        RECT 68.130 3.970 68.550 4.310 ;
        RECT 68.810 4.270 68.980 5.140 ;
        RECT 69.360 4.270 69.530 4.960 ;
        RECT 73.500 4.920 73.670 5.610 ;
        RECT 74.040 4.750 74.210 5.620 ;
        RECT 74.480 5.580 74.900 5.860 ;
        RECT 76.120 5.750 76.290 6.080 ;
        RECT 77.740 5.790 78.000 5.880 ;
        RECT 78.650 5.790 78.910 5.880 ;
        RECT 75.420 5.580 76.840 5.750 ;
        RECT 77.650 5.580 78.070 5.790 ;
        RECT 78.580 5.580 79.000 5.790 ;
        RECT 74.480 5.140 76.060 5.310 ;
        RECT 77.270 5.190 77.440 5.520 ;
        RECT 71.310 4.370 71.480 4.700 ;
        RECT 72.720 4.580 74.300 4.750 ;
        RECT 69.780 4.100 70.200 4.310 ;
        RECT 70.670 4.100 71.090 4.310 ;
        RECT 71.900 4.140 73.360 4.310 ;
        RECT 69.850 4.040 70.110 4.100 ;
        RECT 70.760 4.040 71.020 4.100 ;
        RECT 72.360 4.080 72.650 4.140 ;
        RECT 73.880 3.970 74.300 4.310 ;
        RECT 74.560 4.270 74.730 5.140 ;
        RECT 75.110 4.270 75.280 4.960 ;
        RECT 79.250 4.920 79.420 5.610 ;
        RECT 79.790 4.750 79.960 5.620 ;
        RECT 80.230 5.580 80.650 5.860 ;
        RECT 81.870 5.750 82.040 6.080 ;
        RECT 83.490 5.790 83.750 5.880 ;
        RECT 84.400 5.790 84.660 5.880 ;
        RECT 81.170 5.580 82.590 5.750 ;
        RECT 83.400 5.580 83.820 5.790 ;
        RECT 84.330 5.580 84.750 5.790 ;
        RECT 80.230 5.140 81.810 5.310 ;
        RECT 83.020 5.190 83.190 5.520 ;
        RECT 77.060 4.370 77.230 4.700 ;
        RECT 78.470 4.580 80.050 4.750 ;
        RECT 75.530 4.100 75.950 4.310 ;
        RECT 76.420 4.100 76.840 4.310 ;
        RECT 77.650 4.140 79.110 4.310 ;
        RECT 75.600 4.040 75.860 4.100 ;
        RECT 76.510 4.040 76.770 4.100 ;
        RECT 78.110 4.080 78.400 4.140 ;
        RECT 79.630 3.970 80.050 4.310 ;
        RECT 80.310 4.270 80.480 5.140 ;
        RECT 80.860 4.270 81.030 4.960 ;
        RECT 85.000 4.920 85.170 5.610 ;
        RECT 85.540 4.750 85.710 5.620 ;
        RECT 85.980 5.580 86.400 5.860 ;
        RECT 87.620 5.750 87.790 6.080 ;
        RECT 89.240 5.790 89.500 5.880 ;
        RECT 90.150 5.790 90.410 5.880 ;
        RECT 86.920 5.580 88.340 5.750 ;
        RECT 89.150 5.580 89.570 5.790 ;
        RECT 90.080 5.580 90.500 5.790 ;
        RECT 85.980 5.140 87.560 5.310 ;
        RECT 88.770 5.190 88.940 5.520 ;
        RECT 82.810 4.370 82.980 4.700 ;
        RECT 84.220 4.580 85.800 4.750 ;
        RECT 81.280 4.100 81.700 4.310 ;
        RECT 82.170 4.100 82.590 4.310 ;
        RECT 83.400 4.140 84.860 4.310 ;
        RECT 81.350 4.040 81.610 4.100 ;
        RECT 82.260 4.040 82.520 4.100 ;
        RECT 83.860 4.080 84.150 4.140 ;
        RECT 85.380 3.970 85.800 4.310 ;
        RECT 86.060 4.270 86.230 5.140 ;
        RECT 86.610 4.270 86.780 4.960 ;
        RECT 90.750 4.920 90.920 5.610 ;
        RECT 91.290 4.750 91.460 5.620 ;
        RECT 91.730 5.580 92.150 5.860 ;
        RECT 93.370 5.750 93.540 6.080 ;
        RECT 92.670 5.580 94.090 5.750 ;
        RECT 91.730 5.140 93.310 5.310 ;
        RECT 88.560 4.370 88.730 4.700 ;
        RECT 89.970 4.580 91.550 4.750 ;
        RECT 87.030 4.100 87.450 4.310 ;
        RECT 87.920 4.100 88.340 4.310 ;
        RECT 89.150 4.140 90.610 4.310 ;
        RECT 87.100 4.040 87.360 4.100 ;
        RECT 88.010 4.040 88.270 4.100 ;
        RECT 89.610 4.080 89.900 4.140 ;
        RECT 91.130 3.970 91.550 4.310 ;
        RECT 91.810 4.270 91.980 5.140 ;
        RECT 92.360 4.270 92.530 4.960 ;
        RECT 94.310 4.370 94.480 4.700 ;
        RECT 92.780 4.100 93.200 4.310 ;
        RECT 93.670 4.100 94.090 4.310 ;
        RECT 92.850 4.040 93.110 4.100 ;
        RECT 93.760 4.040 94.020 4.100 ;
        RECT 2.990 3.380 3.250 3.470 ;
        RECT 3.900 3.380 4.160 3.470 ;
        RECT 2.900 3.170 3.320 3.380 ;
        RECT 3.830 3.170 4.250 3.380 ;
        RECT 2.520 2.780 2.690 3.110 ;
        RECT 4.500 2.510 4.670 3.200 ;
        RECT 5.040 2.340 5.210 3.210 ;
        RECT 5.480 3.170 5.900 3.450 ;
        RECT 7.120 3.340 7.290 3.670 ;
        RECT 8.740 3.380 9.000 3.470 ;
        RECT 9.650 3.380 9.910 3.470 ;
        RECT 6.420 3.170 7.840 3.340 ;
        RECT 8.650 3.170 9.070 3.380 ;
        RECT 9.580 3.170 10.000 3.380 ;
        RECT 5.480 2.730 7.060 2.900 ;
        RECT 8.270 2.780 8.440 3.110 ;
        RECT 3.720 2.170 5.300 2.340 ;
        RECT 2.900 1.730 4.360 1.900 ;
        RECT 3.360 1.670 3.650 1.730 ;
        RECT 4.880 1.560 5.300 1.900 ;
        RECT 5.560 1.860 5.730 2.730 ;
        RECT 6.110 1.860 6.280 2.550 ;
        RECT 10.250 2.510 10.420 3.200 ;
        RECT 10.790 2.340 10.960 3.210 ;
        RECT 11.230 3.170 11.650 3.450 ;
        RECT 12.870 3.340 13.040 3.670 ;
        RECT 14.490 3.380 14.750 3.470 ;
        RECT 15.400 3.380 15.660 3.470 ;
        RECT 12.170 3.170 13.590 3.340 ;
        RECT 14.400 3.170 14.820 3.380 ;
        RECT 15.330 3.170 15.750 3.380 ;
        RECT 11.230 2.730 12.810 2.900 ;
        RECT 14.020 2.780 14.190 3.110 ;
        RECT 8.060 1.960 8.230 2.290 ;
        RECT 9.470 2.170 11.050 2.340 ;
        RECT 6.530 1.690 6.950 1.900 ;
        RECT 7.420 1.690 7.840 1.900 ;
        RECT 8.650 1.730 10.110 1.900 ;
        RECT 6.600 1.630 6.860 1.690 ;
        RECT 7.510 1.630 7.770 1.690 ;
        RECT 9.110 1.670 9.400 1.730 ;
        RECT 10.630 1.560 11.050 1.900 ;
        RECT 11.310 1.860 11.480 2.730 ;
        RECT 11.860 1.860 12.030 2.550 ;
        RECT 16.000 2.510 16.170 3.200 ;
        RECT 16.540 2.340 16.710 3.210 ;
        RECT 16.980 3.170 17.400 3.450 ;
        RECT 18.620 3.340 18.790 3.670 ;
        RECT 20.240 3.380 20.500 3.470 ;
        RECT 21.150 3.380 21.410 3.470 ;
        RECT 17.920 3.170 19.340 3.340 ;
        RECT 20.150 3.170 20.570 3.380 ;
        RECT 21.080 3.170 21.500 3.380 ;
        RECT 16.980 2.730 18.560 2.900 ;
        RECT 19.770 2.780 19.940 3.110 ;
        RECT 13.810 1.960 13.980 2.290 ;
        RECT 15.220 2.170 16.800 2.340 ;
        RECT 12.280 1.690 12.700 1.900 ;
        RECT 13.170 1.690 13.590 1.900 ;
        RECT 14.400 1.730 15.860 1.900 ;
        RECT 12.350 1.630 12.610 1.690 ;
        RECT 13.260 1.630 13.520 1.690 ;
        RECT 14.860 1.670 15.150 1.730 ;
        RECT 16.380 1.560 16.800 1.900 ;
        RECT 17.060 1.860 17.230 2.730 ;
        RECT 17.610 1.860 17.780 2.550 ;
        RECT 21.750 2.510 21.920 3.200 ;
        RECT 22.290 2.340 22.460 3.210 ;
        RECT 22.730 3.170 23.150 3.450 ;
        RECT 24.370 3.340 24.540 3.670 ;
        RECT 25.990 3.380 26.250 3.470 ;
        RECT 26.900 3.380 27.160 3.470 ;
        RECT 23.670 3.170 25.090 3.340 ;
        RECT 25.900 3.170 26.320 3.380 ;
        RECT 26.830 3.170 27.250 3.380 ;
        RECT 22.730 2.730 24.310 2.900 ;
        RECT 25.520 2.780 25.690 3.110 ;
        RECT 19.560 1.960 19.730 2.290 ;
        RECT 20.970 2.170 22.550 2.340 ;
        RECT 18.030 1.690 18.450 1.900 ;
        RECT 18.920 1.690 19.340 1.900 ;
        RECT 20.150 1.730 21.610 1.900 ;
        RECT 18.100 1.630 18.360 1.690 ;
        RECT 19.010 1.630 19.270 1.690 ;
        RECT 20.610 1.670 20.900 1.730 ;
        RECT 22.130 1.560 22.550 1.900 ;
        RECT 22.810 1.860 22.980 2.730 ;
        RECT 23.360 1.860 23.530 2.550 ;
        RECT 27.500 2.510 27.670 3.200 ;
        RECT 28.040 2.340 28.210 3.210 ;
        RECT 28.480 3.170 28.900 3.450 ;
        RECT 30.120 3.340 30.290 3.670 ;
        RECT 31.740 3.380 32.000 3.470 ;
        RECT 32.650 3.380 32.910 3.470 ;
        RECT 29.420 3.170 30.840 3.340 ;
        RECT 31.650 3.170 32.070 3.380 ;
        RECT 32.580 3.170 33.000 3.380 ;
        RECT 28.480 2.730 30.060 2.900 ;
        RECT 31.270 2.780 31.440 3.110 ;
        RECT 25.310 1.960 25.480 2.290 ;
        RECT 26.720 2.170 28.300 2.340 ;
        RECT 23.780 1.690 24.200 1.900 ;
        RECT 24.670 1.690 25.090 1.900 ;
        RECT 25.900 1.730 27.360 1.900 ;
        RECT 23.850 1.630 24.110 1.690 ;
        RECT 24.760 1.630 25.020 1.690 ;
        RECT 26.360 1.670 26.650 1.730 ;
        RECT 27.880 1.560 28.300 1.900 ;
        RECT 28.560 1.860 28.730 2.730 ;
        RECT 29.110 1.860 29.280 2.550 ;
        RECT 33.250 2.510 33.420 3.200 ;
        RECT 33.790 2.340 33.960 3.210 ;
        RECT 34.230 3.170 34.650 3.450 ;
        RECT 35.870 3.340 36.040 3.670 ;
        RECT 37.490 3.380 37.750 3.470 ;
        RECT 38.400 3.380 38.660 3.470 ;
        RECT 35.170 3.170 36.590 3.340 ;
        RECT 37.400 3.170 37.820 3.380 ;
        RECT 38.330 3.170 38.750 3.380 ;
        RECT 34.230 2.730 35.810 2.900 ;
        RECT 37.020 2.780 37.190 3.110 ;
        RECT 31.060 1.960 31.230 2.290 ;
        RECT 32.470 2.170 34.050 2.340 ;
        RECT 29.530 1.690 29.950 1.900 ;
        RECT 30.420 1.690 30.840 1.900 ;
        RECT 31.650 1.730 33.110 1.900 ;
        RECT 29.600 1.630 29.860 1.690 ;
        RECT 30.510 1.630 30.770 1.690 ;
        RECT 32.110 1.670 32.400 1.730 ;
        RECT 33.630 1.560 34.050 1.900 ;
        RECT 34.310 1.860 34.480 2.730 ;
        RECT 34.860 1.860 35.030 2.550 ;
        RECT 39.000 2.510 39.170 3.200 ;
        RECT 39.540 2.340 39.710 3.210 ;
        RECT 39.980 3.170 40.400 3.450 ;
        RECT 41.620 3.340 41.790 3.670 ;
        RECT 43.240 3.380 43.500 3.470 ;
        RECT 44.150 3.380 44.410 3.470 ;
        RECT 40.920 3.170 42.340 3.340 ;
        RECT 43.150 3.170 43.570 3.380 ;
        RECT 44.080 3.170 44.500 3.380 ;
        RECT 39.980 2.730 41.560 2.900 ;
        RECT 42.770 2.780 42.940 3.110 ;
        RECT 36.810 1.960 36.980 2.290 ;
        RECT 38.220 2.170 39.800 2.340 ;
        RECT 35.280 1.690 35.700 1.900 ;
        RECT 36.170 1.690 36.590 1.900 ;
        RECT 37.400 1.730 38.860 1.900 ;
        RECT 35.350 1.630 35.610 1.690 ;
        RECT 36.260 1.630 36.520 1.690 ;
        RECT 37.860 1.670 38.150 1.730 ;
        RECT 39.380 1.560 39.800 1.900 ;
        RECT 40.060 1.860 40.230 2.730 ;
        RECT 40.610 1.860 40.780 2.550 ;
        RECT 44.750 2.510 44.920 3.200 ;
        RECT 45.290 2.340 45.460 3.210 ;
        RECT 45.730 3.170 46.150 3.450 ;
        RECT 47.370 3.340 47.540 3.670 ;
        RECT 48.990 3.380 49.250 3.470 ;
        RECT 49.900 3.380 50.160 3.470 ;
        RECT 46.670 3.170 48.090 3.340 ;
        RECT 48.900 3.170 49.320 3.380 ;
        RECT 49.830 3.170 50.250 3.380 ;
        RECT 45.730 2.730 47.310 2.900 ;
        RECT 48.520 2.780 48.690 3.110 ;
        RECT 42.560 1.960 42.730 2.290 ;
        RECT 43.970 2.170 45.550 2.340 ;
        RECT 41.030 1.690 41.450 1.900 ;
        RECT 41.920 1.690 42.340 1.900 ;
        RECT 43.150 1.730 44.610 1.900 ;
        RECT 41.100 1.630 41.360 1.690 ;
        RECT 42.010 1.630 42.270 1.690 ;
        RECT 43.610 1.670 43.900 1.730 ;
        RECT 45.130 1.560 45.550 1.900 ;
        RECT 45.810 1.860 45.980 2.730 ;
        RECT 46.360 1.860 46.530 2.550 ;
        RECT 50.500 2.510 50.670 3.200 ;
        RECT 51.040 2.340 51.210 3.210 ;
        RECT 51.480 3.170 51.900 3.450 ;
        RECT 53.120 3.340 53.290 3.670 ;
        RECT 54.740 3.380 55.000 3.470 ;
        RECT 55.650 3.380 55.910 3.470 ;
        RECT 52.420 3.170 53.840 3.340 ;
        RECT 54.650 3.170 55.070 3.380 ;
        RECT 55.580 3.170 56.000 3.380 ;
        RECT 51.480 2.730 53.060 2.900 ;
        RECT 54.270 2.780 54.440 3.110 ;
        RECT 48.310 1.960 48.480 2.290 ;
        RECT 49.720 2.170 51.300 2.340 ;
        RECT 46.780 1.690 47.200 1.900 ;
        RECT 47.670 1.690 48.090 1.900 ;
        RECT 48.900 1.730 50.360 1.900 ;
        RECT 46.850 1.630 47.110 1.690 ;
        RECT 47.760 1.630 48.020 1.690 ;
        RECT 49.360 1.670 49.650 1.730 ;
        RECT 50.880 1.560 51.300 1.900 ;
        RECT 51.560 1.860 51.730 2.730 ;
        RECT 52.110 1.860 52.280 2.550 ;
        RECT 56.250 2.510 56.420 3.200 ;
        RECT 56.790 2.340 56.960 3.210 ;
        RECT 57.230 3.170 57.650 3.450 ;
        RECT 58.870 3.340 59.040 3.670 ;
        RECT 60.490 3.380 60.750 3.470 ;
        RECT 61.400 3.380 61.660 3.470 ;
        RECT 58.170 3.170 59.590 3.340 ;
        RECT 60.400 3.170 60.820 3.380 ;
        RECT 61.330 3.170 61.750 3.380 ;
        RECT 57.230 2.730 58.810 2.900 ;
        RECT 60.020 2.780 60.190 3.110 ;
        RECT 54.060 1.960 54.230 2.290 ;
        RECT 55.470 2.170 57.050 2.340 ;
        RECT 52.530 1.690 52.950 1.900 ;
        RECT 53.420 1.690 53.840 1.900 ;
        RECT 54.650 1.730 56.110 1.900 ;
        RECT 52.600 1.630 52.860 1.690 ;
        RECT 53.510 1.630 53.770 1.690 ;
        RECT 55.110 1.670 55.400 1.730 ;
        RECT 56.630 1.560 57.050 1.900 ;
        RECT 57.310 1.860 57.480 2.730 ;
        RECT 57.860 1.860 58.030 2.550 ;
        RECT 62.000 2.510 62.170 3.200 ;
        RECT 62.540 2.340 62.710 3.210 ;
        RECT 62.980 3.170 63.400 3.450 ;
        RECT 64.620 3.340 64.790 3.670 ;
        RECT 66.240 3.380 66.500 3.470 ;
        RECT 67.150 3.380 67.410 3.470 ;
        RECT 63.920 3.170 65.340 3.340 ;
        RECT 66.150 3.170 66.570 3.380 ;
        RECT 67.080 3.170 67.500 3.380 ;
        RECT 62.980 2.730 64.560 2.900 ;
        RECT 65.770 2.780 65.940 3.110 ;
        RECT 59.810 1.960 59.980 2.290 ;
        RECT 61.220 2.170 62.800 2.340 ;
        RECT 58.280 1.690 58.700 1.900 ;
        RECT 59.170 1.690 59.590 1.900 ;
        RECT 60.400 1.730 61.860 1.900 ;
        RECT 58.350 1.630 58.610 1.690 ;
        RECT 59.260 1.630 59.520 1.690 ;
        RECT 60.860 1.670 61.150 1.730 ;
        RECT 62.380 1.560 62.800 1.900 ;
        RECT 63.060 1.860 63.230 2.730 ;
        RECT 63.610 1.860 63.780 2.550 ;
        RECT 67.750 2.510 67.920 3.200 ;
        RECT 68.290 2.340 68.460 3.210 ;
        RECT 68.730 3.170 69.150 3.450 ;
        RECT 70.370 3.340 70.540 3.670 ;
        RECT 71.990 3.380 72.250 3.470 ;
        RECT 72.900 3.380 73.160 3.470 ;
        RECT 69.670 3.170 71.090 3.340 ;
        RECT 71.900 3.170 72.320 3.380 ;
        RECT 72.830 3.170 73.250 3.380 ;
        RECT 68.730 2.730 70.310 2.900 ;
        RECT 71.520 2.780 71.690 3.110 ;
        RECT 65.560 1.960 65.730 2.290 ;
        RECT 66.970 2.170 68.550 2.340 ;
        RECT 64.030 1.690 64.450 1.900 ;
        RECT 64.920 1.690 65.340 1.900 ;
        RECT 66.150 1.730 67.610 1.900 ;
        RECT 64.100 1.630 64.360 1.690 ;
        RECT 65.010 1.630 65.270 1.690 ;
        RECT 66.610 1.670 66.900 1.730 ;
        RECT 68.130 1.560 68.550 1.900 ;
        RECT 68.810 1.860 68.980 2.730 ;
        RECT 69.360 1.860 69.530 2.550 ;
        RECT 73.500 2.510 73.670 3.200 ;
        RECT 74.040 2.340 74.210 3.210 ;
        RECT 74.480 3.170 74.900 3.450 ;
        RECT 76.120 3.340 76.290 3.670 ;
        RECT 77.740 3.380 78.000 3.470 ;
        RECT 78.650 3.380 78.910 3.470 ;
        RECT 75.420 3.170 76.840 3.340 ;
        RECT 77.650 3.170 78.070 3.380 ;
        RECT 78.580 3.170 79.000 3.380 ;
        RECT 74.480 2.730 76.060 2.900 ;
        RECT 77.270 2.780 77.440 3.110 ;
        RECT 71.310 1.960 71.480 2.290 ;
        RECT 72.720 2.170 74.300 2.340 ;
        RECT 69.780 1.690 70.200 1.900 ;
        RECT 70.670 1.690 71.090 1.900 ;
        RECT 71.900 1.730 73.360 1.900 ;
        RECT 69.850 1.630 70.110 1.690 ;
        RECT 70.760 1.630 71.020 1.690 ;
        RECT 72.360 1.670 72.650 1.730 ;
        RECT 73.880 1.560 74.300 1.900 ;
        RECT 74.560 1.860 74.730 2.730 ;
        RECT 75.110 1.860 75.280 2.550 ;
        RECT 79.250 2.510 79.420 3.200 ;
        RECT 79.790 2.340 79.960 3.210 ;
        RECT 80.230 3.170 80.650 3.450 ;
        RECT 81.870 3.340 82.040 3.670 ;
        RECT 83.490 3.380 83.750 3.470 ;
        RECT 84.400 3.380 84.660 3.470 ;
        RECT 81.170 3.170 82.590 3.340 ;
        RECT 83.400 3.170 83.820 3.380 ;
        RECT 84.330 3.170 84.750 3.380 ;
        RECT 80.230 2.730 81.810 2.900 ;
        RECT 83.020 2.780 83.190 3.110 ;
        RECT 77.060 1.960 77.230 2.290 ;
        RECT 78.470 2.170 80.050 2.340 ;
        RECT 75.530 1.690 75.950 1.900 ;
        RECT 76.420 1.690 76.840 1.900 ;
        RECT 77.650 1.730 79.110 1.900 ;
        RECT 75.600 1.630 75.860 1.690 ;
        RECT 76.510 1.630 76.770 1.690 ;
        RECT 78.110 1.670 78.400 1.730 ;
        RECT 79.630 1.560 80.050 1.900 ;
        RECT 80.310 1.860 80.480 2.730 ;
        RECT 80.860 1.860 81.030 2.550 ;
        RECT 85.000 2.510 85.170 3.200 ;
        RECT 85.540 2.340 85.710 3.210 ;
        RECT 85.980 3.170 86.400 3.450 ;
        RECT 87.620 3.340 87.790 3.670 ;
        RECT 89.240 3.380 89.500 3.470 ;
        RECT 90.150 3.380 90.410 3.470 ;
        RECT 86.920 3.170 88.340 3.340 ;
        RECT 89.150 3.170 89.570 3.380 ;
        RECT 90.080 3.170 90.500 3.380 ;
        RECT 85.980 2.730 87.560 2.900 ;
        RECT 88.770 2.780 88.940 3.110 ;
        RECT 82.810 1.960 82.980 2.290 ;
        RECT 84.220 2.170 85.800 2.340 ;
        RECT 81.280 1.690 81.700 1.900 ;
        RECT 82.170 1.690 82.590 1.900 ;
        RECT 83.400 1.730 84.860 1.900 ;
        RECT 81.350 1.630 81.610 1.690 ;
        RECT 82.260 1.630 82.520 1.690 ;
        RECT 83.860 1.670 84.150 1.730 ;
        RECT 85.380 1.560 85.800 1.900 ;
        RECT 86.060 1.860 86.230 2.730 ;
        RECT 86.610 1.860 86.780 2.550 ;
        RECT 90.750 2.510 90.920 3.200 ;
        RECT 91.290 2.340 91.460 3.210 ;
        RECT 91.730 3.170 92.150 3.450 ;
        RECT 93.370 3.340 93.540 3.670 ;
        RECT 92.670 3.170 94.090 3.340 ;
        RECT 91.730 2.730 93.310 2.900 ;
        RECT 88.560 1.960 88.730 2.290 ;
        RECT 89.970 2.170 91.550 2.340 ;
        RECT 87.030 1.690 87.450 1.900 ;
        RECT 87.920 1.690 88.340 1.900 ;
        RECT 89.150 1.730 90.610 1.900 ;
        RECT 87.100 1.630 87.360 1.690 ;
        RECT 88.010 1.630 88.270 1.690 ;
        RECT 89.610 1.670 89.900 1.730 ;
        RECT 91.130 1.560 91.550 1.900 ;
        RECT 91.810 1.860 91.980 2.730 ;
        RECT 92.360 1.860 92.530 2.550 ;
        RECT 94.310 1.960 94.480 2.290 ;
        RECT 92.780 1.690 93.200 1.900 ;
        RECT 93.670 1.690 94.090 1.900 ;
        RECT 92.850 1.630 93.110 1.690 ;
        RECT 93.760 1.630 94.020 1.690 ;
        RECT 2.990 0.970 3.250 1.060 ;
        RECT 3.900 0.970 4.160 1.060 ;
        RECT 2.900 0.760 3.320 0.970 ;
        RECT 3.830 0.760 4.250 0.970 ;
        RECT 2.520 0.370 2.690 0.700 ;
        RECT 4.500 0.100 4.670 0.790 ;
        RECT 5.040 -0.070 5.210 0.800 ;
        RECT 5.480 0.760 5.900 1.040 ;
        RECT 7.120 0.930 7.290 1.260 ;
        RECT 8.740 0.970 9.000 1.060 ;
        RECT 9.650 0.970 9.910 1.060 ;
        RECT 6.420 0.760 7.840 0.930 ;
        RECT 8.650 0.760 9.070 0.970 ;
        RECT 9.580 0.760 10.000 0.970 ;
        RECT 5.480 0.320 7.060 0.490 ;
        RECT 8.270 0.370 8.440 0.700 ;
        RECT 3.720 -0.240 5.300 -0.070 ;
        RECT 2.900 -0.680 4.360 -0.510 ;
        RECT 3.360 -0.740 3.650 -0.680 ;
        RECT 4.880 -0.850 5.300 -0.510 ;
        RECT 5.560 -0.550 5.730 0.320 ;
        RECT 6.110 -0.550 6.280 0.140 ;
        RECT 10.250 0.100 10.420 0.790 ;
        RECT 10.790 -0.070 10.960 0.800 ;
        RECT 11.230 0.760 11.650 1.040 ;
        RECT 12.870 0.930 13.040 1.260 ;
        RECT 14.490 0.970 14.750 1.060 ;
        RECT 15.400 0.970 15.660 1.060 ;
        RECT 12.170 0.760 13.590 0.930 ;
        RECT 14.400 0.760 14.820 0.970 ;
        RECT 15.330 0.760 15.750 0.970 ;
        RECT 11.230 0.320 12.810 0.490 ;
        RECT 14.020 0.370 14.190 0.700 ;
        RECT 8.060 -0.450 8.230 -0.120 ;
        RECT 9.470 -0.240 11.050 -0.070 ;
        RECT 6.530 -0.720 6.950 -0.510 ;
        RECT 7.420 -0.720 7.840 -0.510 ;
        RECT 8.650 -0.680 10.110 -0.510 ;
        RECT 6.600 -0.780 6.860 -0.720 ;
        RECT 7.510 -0.780 7.770 -0.720 ;
        RECT 9.110 -0.740 9.400 -0.680 ;
        RECT 10.630 -0.850 11.050 -0.510 ;
        RECT 11.310 -0.550 11.480 0.320 ;
        RECT 11.860 -0.550 12.030 0.140 ;
        RECT 16.000 0.100 16.170 0.790 ;
        RECT 16.540 -0.070 16.710 0.800 ;
        RECT 16.980 0.760 17.400 1.040 ;
        RECT 18.620 0.930 18.790 1.260 ;
        RECT 20.240 0.970 20.500 1.060 ;
        RECT 21.150 0.970 21.410 1.060 ;
        RECT 17.920 0.760 19.340 0.930 ;
        RECT 20.150 0.760 20.570 0.970 ;
        RECT 21.080 0.760 21.500 0.970 ;
        RECT 16.980 0.320 18.560 0.490 ;
        RECT 19.770 0.370 19.940 0.700 ;
        RECT 13.810 -0.450 13.980 -0.120 ;
        RECT 15.220 -0.240 16.800 -0.070 ;
        RECT 12.280 -0.720 12.700 -0.510 ;
        RECT 13.170 -0.720 13.590 -0.510 ;
        RECT 14.400 -0.680 15.860 -0.510 ;
        RECT 12.350 -0.780 12.610 -0.720 ;
        RECT 13.260 -0.780 13.520 -0.720 ;
        RECT 14.860 -0.740 15.150 -0.680 ;
        RECT 16.380 -0.850 16.800 -0.510 ;
        RECT 17.060 -0.550 17.230 0.320 ;
        RECT 17.610 -0.550 17.780 0.140 ;
        RECT 21.750 0.100 21.920 0.790 ;
        RECT 22.290 -0.070 22.460 0.800 ;
        RECT 22.730 0.760 23.150 1.040 ;
        RECT 24.370 0.930 24.540 1.260 ;
        RECT 25.990 0.970 26.250 1.060 ;
        RECT 26.900 0.970 27.160 1.060 ;
        RECT 23.670 0.760 25.090 0.930 ;
        RECT 25.900 0.760 26.320 0.970 ;
        RECT 26.830 0.760 27.250 0.970 ;
        RECT 22.730 0.320 24.310 0.490 ;
        RECT 25.520 0.370 25.690 0.700 ;
        RECT 19.560 -0.450 19.730 -0.120 ;
        RECT 20.970 -0.240 22.550 -0.070 ;
        RECT 18.030 -0.720 18.450 -0.510 ;
        RECT 18.920 -0.720 19.340 -0.510 ;
        RECT 20.150 -0.680 21.610 -0.510 ;
        RECT 18.100 -0.780 18.360 -0.720 ;
        RECT 19.010 -0.780 19.270 -0.720 ;
        RECT 20.610 -0.740 20.900 -0.680 ;
        RECT 22.130 -0.850 22.550 -0.510 ;
        RECT 22.810 -0.550 22.980 0.320 ;
        RECT 23.360 -0.550 23.530 0.140 ;
        RECT 27.500 0.100 27.670 0.790 ;
        RECT 28.040 -0.070 28.210 0.800 ;
        RECT 28.480 0.760 28.900 1.040 ;
        RECT 30.120 0.930 30.290 1.260 ;
        RECT 31.740 0.970 32.000 1.060 ;
        RECT 32.650 0.970 32.910 1.060 ;
        RECT 29.420 0.760 30.840 0.930 ;
        RECT 31.650 0.760 32.070 0.970 ;
        RECT 32.580 0.760 33.000 0.970 ;
        RECT 28.480 0.320 30.060 0.490 ;
        RECT 31.270 0.370 31.440 0.700 ;
        RECT 25.310 -0.450 25.480 -0.120 ;
        RECT 26.720 -0.240 28.300 -0.070 ;
        RECT 23.780 -0.720 24.200 -0.510 ;
        RECT 24.670 -0.720 25.090 -0.510 ;
        RECT 25.900 -0.680 27.360 -0.510 ;
        RECT 23.850 -0.780 24.110 -0.720 ;
        RECT 24.760 -0.780 25.020 -0.720 ;
        RECT 26.360 -0.740 26.650 -0.680 ;
        RECT 27.880 -0.850 28.300 -0.510 ;
        RECT 28.560 -0.550 28.730 0.320 ;
        RECT 29.110 -0.550 29.280 0.140 ;
        RECT 33.250 0.100 33.420 0.790 ;
        RECT 33.790 -0.070 33.960 0.800 ;
        RECT 34.230 0.760 34.650 1.040 ;
        RECT 35.870 0.930 36.040 1.260 ;
        RECT 37.490 0.970 37.750 1.060 ;
        RECT 38.400 0.970 38.660 1.060 ;
        RECT 35.170 0.760 36.590 0.930 ;
        RECT 37.400 0.760 37.820 0.970 ;
        RECT 38.330 0.760 38.750 0.970 ;
        RECT 34.230 0.320 35.810 0.490 ;
        RECT 37.020 0.370 37.190 0.700 ;
        RECT 31.060 -0.450 31.230 -0.120 ;
        RECT 32.470 -0.240 34.050 -0.070 ;
        RECT 29.530 -0.720 29.950 -0.510 ;
        RECT 30.420 -0.720 30.840 -0.510 ;
        RECT 31.650 -0.680 33.110 -0.510 ;
        RECT 29.600 -0.780 29.860 -0.720 ;
        RECT 30.510 -0.780 30.770 -0.720 ;
        RECT 32.110 -0.740 32.400 -0.680 ;
        RECT 33.630 -0.850 34.050 -0.510 ;
        RECT 34.310 -0.550 34.480 0.320 ;
        RECT 34.860 -0.550 35.030 0.140 ;
        RECT 39.000 0.100 39.170 0.790 ;
        RECT 39.540 -0.070 39.710 0.800 ;
        RECT 39.980 0.760 40.400 1.040 ;
        RECT 41.620 0.930 41.790 1.260 ;
        RECT 43.240 0.970 43.500 1.060 ;
        RECT 44.150 0.970 44.410 1.060 ;
        RECT 40.920 0.760 42.340 0.930 ;
        RECT 43.150 0.760 43.570 0.970 ;
        RECT 44.080 0.760 44.500 0.970 ;
        RECT 39.980 0.320 41.560 0.490 ;
        RECT 42.770 0.370 42.940 0.700 ;
        RECT 36.810 -0.450 36.980 -0.120 ;
        RECT 38.220 -0.240 39.800 -0.070 ;
        RECT 35.280 -0.720 35.700 -0.510 ;
        RECT 36.170 -0.720 36.590 -0.510 ;
        RECT 37.400 -0.680 38.860 -0.510 ;
        RECT 35.350 -0.780 35.610 -0.720 ;
        RECT 36.260 -0.780 36.520 -0.720 ;
        RECT 37.860 -0.740 38.150 -0.680 ;
        RECT 39.380 -0.850 39.800 -0.510 ;
        RECT 40.060 -0.550 40.230 0.320 ;
        RECT 40.610 -0.550 40.780 0.140 ;
        RECT 44.750 0.100 44.920 0.790 ;
        RECT 45.290 -0.070 45.460 0.800 ;
        RECT 45.730 0.760 46.150 1.040 ;
        RECT 47.370 0.930 47.540 1.260 ;
        RECT 48.990 0.970 49.250 1.060 ;
        RECT 49.900 0.970 50.160 1.060 ;
        RECT 46.670 0.760 48.090 0.930 ;
        RECT 48.900 0.760 49.320 0.970 ;
        RECT 49.830 0.760 50.250 0.970 ;
        RECT 45.730 0.320 47.310 0.490 ;
        RECT 48.520 0.370 48.690 0.700 ;
        RECT 42.560 -0.450 42.730 -0.120 ;
        RECT 43.970 -0.240 45.550 -0.070 ;
        RECT 41.030 -0.720 41.450 -0.510 ;
        RECT 41.920 -0.720 42.340 -0.510 ;
        RECT 43.150 -0.680 44.610 -0.510 ;
        RECT 41.100 -0.780 41.360 -0.720 ;
        RECT 42.010 -0.780 42.270 -0.720 ;
        RECT 43.610 -0.740 43.900 -0.680 ;
        RECT 45.130 -0.850 45.550 -0.510 ;
        RECT 45.810 -0.550 45.980 0.320 ;
        RECT 46.360 -0.550 46.530 0.140 ;
        RECT 50.500 0.100 50.670 0.790 ;
        RECT 51.040 -0.070 51.210 0.800 ;
        RECT 51.480 0.760 51.900 1.040 ;
        RECT 53.120 0.930 53.290 1.260 ;
        RECT 54.740 0.970 55.000 1.060 ;
        RECT 55.650 0.970 55.910 1.060 ;
        RECT 52.420 0.760 53.840 0.930 ;
        RECT 54.650 0.760 55.070 0.970 ;
        RECT 55.580 0.760 56.000 0.970 ;
        RECT 51.480 0.320 53.060 0.490 ;
        RECT 54.270 0.370 54.440 0.700 ;
        RECT 48.310 -0.450 48.480 -0.120 ;
        RECT 49.720 -0.240 51.300 -0.070 ;
        RECT 46.780 -0.720 47.200 -0.510 ;
        RECT 47.670 -0.720 48.090 -0.510 ;
        RECT 48.900 -0.680 50.360 -0.510 ;
        RECT 46.850 -0.780 47.110 -0.720 ;
        RECT 47.760 -0.780 48.020 -0.720 ;
        RECT 49.360 -0.740 49.650 -0.680 ;
        RECT 50.880 -0.850 51.300 -0.510 ;
        RECT 51.560 -0.550 51.730 0.320 ;
        RECT 52.110 -0.550 52.280 0.140 ;
        RECT 56.250 0.100 56.420 0.790 ;
        RECT 56.790 -0.070 56.960 0.800 ;
        RECT 57.230 0.760 57.650 1.040 ;
        RECT 58.870 0.930 59.040 1.260 ;
        RECT 60.490 0.970 60.750 1.060 ;
        RECT 61.400 0.970 61.660 1.060 ;
        RECT 58.170 0.760 59.590 0.930 ;
        RECT 60.400 0.760 60.820 0.970 ;
        RECT 61.330 0.760 61.750 0.970 ;
        RECT 57.230 0.320 58.810 0.490 ;
        RECT 60.020 0.370 60.190 0.700 ;
        RECT 54.060 -0.450 54.230 -0.120 ;
        RECT 55.470 -0.240 57.050 -0.070 ;
        RECT 52.530 -0.720 52.950 -0.510 ;
        RECT 53.420 -0.720 53.840 -0.510 ;
        RECT 54.650 -0.680 56.110 -0.510 ;
        RECT 52.600 -0.780 52.860 -0.720 ;
        RECT 53.510 -0.780 53.770 -0.720 ;
        RECT 55.110 -0.740 55.400 -0.680 ;
        RECT 56.630 -0.850 57.050 -0.510 ;
        RECT 57.310 -0.550 57.480 0.320 ;
        RECT 57.860 -0.550 58.030 0.140 ;
        RECT 62.000 0.100 62.170 0.790 ;
        RECT 62.540 -0.070 62.710 0.800 ;
        RECT 62.980 0.760 63.400 1.040 ;
        RECT 64.620 0.930 64.790 1.260 ;
        RECT 66.240 0.970 66.500 1.060 ;
        RECT 67.150 0.970 67.410 1.060 ;
        RECT 63.920 0.760 65.340 0.930 ;
        RECT 66.150 0.760 66.570 0.970 ;
        RECT 67.080 0.760 67.500 0.970 ;
        RECT 62.980 0.320 64.560 0.490 ;
        RECT 65.770 0.370 65.940 0.700 ;
        RECT 59.810 -0.450 59.980 -0.120 ;
        RECT 61.220 -0.240 62.800 -0.070 ;
        RECT 58.280 -0.720 58.700 -0.510 ;
        RECT 59.170 -0.720 59.590 -0.510 ;
        RECT 60.400 -0.680 61.860 -0.510 ;
        RECT 58.350 -0.780 58.610 -0.720 ;
        RECT 59.260 -0.780 59.520 -0.720 ;
        RECT 60.860 -0.740 61.150 -0.680 ;
        RECT 62.380 -0.850 62.800 -0.510 ;
        RECT 63.060 -0.550 63.230 0.320 ;
        RECT 63.610 -0.550 63.780 0.140 ;
        RECT 67.750 0.100 67.920 0.790 ;
        RECT 68.290 -0.070 68.460 0.800 ;
        RECT 68.730 0.760 69.150 1.040 ;
        RECT 70.370 0.930 70.540 1.260 ;
        RECT 71.990 0.970 72.250 1.060 ;
        RECT 72.900 0.970 73.160 1.060 ;
        RECT 69.670 0.760 71.090 0.930 ;
        RECT 71.900 0.760 72.320 0.970 ;
        RECT 72.830 0.760 73.250 0.970 ;
        RECT 68.730 0.320 70.310 0.490 ;
        RECT 71.520 0.370 71.690 0.700 ;
        RECT 65.560 -0.450 65.730 -0.120 ;
        RECT 66.970 -0.240 68.550 -0.070 ;
        RECT 64.030 -0.720 64.450 -0.510 ;
        RECT 64.920 -0.720 65.340 -0.510 ;
        RECT 66.150 -0.680 67.610 -0.510 ;
        RECT 64.100 -0.780 64.360 -0.720 ;
        RECT 65.010 -0.780 65.270 -0.720 ;
        RECT 66.610 -0.740 66.900 -0.680 ;
        RECT 68.130 -0.850 68.550 -0.510 ;
        RECT 68.810 -0.550 68.980 0.320 ;
        RECT 69.360 -0.550 69.530 0.140 ;
        RECT 73.500 0.100 73.670 0.790 ;
        RECT 74.040 -0.070 74.210 0.800 ;
        RECT 74.480 0.760 74.900 1.040 ;
        RECT 76.120 0.930 76.290 1.260 ;
        RECT 77.740 0.970 78.000 1.060 ;
        RECT 78.650 0.970 78.910 1.060 ;
        RECT 75.420 0.760 76.840 0.930 ;
        RECT 77.650 0.760 78.070 0.970 ;
        RECT 78.580 0.760 79.000 0.970 ;
        RECT 74.480 0.320 76.060 0.490 ;
        RECT 77.270 0.370 77.440 0.700 ;
        RECT 71.310 -0.450 71.480 -0.120 ;
        RECT 72.720 -0.240 74.300 -0.070 ;
        RECT 69.780 -0.720 70.200 -0.510 ;
        RECT 70.670 -0.720 71.090 -0.510 ;
        RECT 71.900 -0.680 73.360 -0.510 ;
        RECT 69.850 -0.780 70.110 -0.720 ;
        RECT 70.760 -0.780 71.020 -0.720 ;
        RECT 72.360 -0.740 72.650 -0.680 ;
        RECT 73.880 -0.850 74.300 -0.510 ;
        RECT 74.560 -0.550 74.730 0.320 ;
        RECT 75.110 -0.550 75.280 0.140 ;
        RECT 79.250 0.100 79.420 0.790 ;
        RECT 79.790 -0.070 79.960 0.800 ;
        RECT 80.230 0.760 80.650 1.040 ;
        RECT 81.870 0.930 82.040 1.260 ;
        RECT 83.490 0.970 83.750 1.060 ;
        RECT 84.400 0.970 84.660 1.060 ;
        RECT 81.170 0.760 82.590 0.930 ;
        RECT 83.400 0.760 83.820 0.970 ;
        RECT 84.330 0.760 84.750 0.970 ;
        RECT 80.230 0.320 81.810 0.490 ;
        RECT 83.020 0.370 83.190 0.700 ;
        RECT 77.060 -0.450 77.230 -0.120 ;
        RECT 78.470 -0.240 80.050 -0.070 ;
        RECT 75.530 -0.720 75.950 -0.510 ;
        RECT 76.420 -0.720 76.840 -0.510 ;
        RECT 77.650 -0.680 79.110 -0.510 ;
        RECT 75.600 -0.780 75.860 -0.720 ;
        RECT 76.510 -0.780 76.770 -0.720 ;
        RECT 78.110 -0.740 78.400 -0.680 ;
        RECT 79.630 -0.850 80.050 -0.510 ;
        RECT 80.310 -0.550 80.480 0.320 ;
        RECT 80.860 -0.550 81.030 0.140 ;
        RECT 85.000 0.100 85.170 0.790 ;
        RECT 85.540 -0.070 85.710 0.800 ;
        RECT 85.980 0.760 86.400 1.040 ;
        RECT 87.620 0.930 87.790 1.260 ;
        RECT 89.240 0.970 89.500 1.060 ;
        RECT 90.150 0.970 90.410 1.060 ;
        RECT 86.920 0.760 88.340 0.930 ;
        RECT 89.150 0.760 89.570 0.970 ;
        RECT 90.080 0.760 90.500 0.970 ;
        RECT 85.980 0.320 87.560 0.490 ;
        RECT 88.770 0.370 88.940 0.700 ;
        RECT 82.810 -0.450 82.980 -0.120 ;
        RECT 84.220 -0.240 85.800 -0.070 ;
        RECT 81.280 -0.720 81.700 -0.510 ;
        RECT 82.170 -0.720 82.590 -0.510 ;
        RECT 83.400 -0.680 84.860 -0.510 ;
        RECT 81.350 -0.780 81.610 -0.720 ;
        RECT 82.260 -0.780 82.520 -0.720 ;
        RECT 83.860 -0.740 84.150 -0.680 ;
        RECT 85.380 -0.850 85.800 -0.510 ;
        RECT 86.060 -0.550 86.230 0.320 ;
        RECT 86.610 -0.550 86.780 0.140 ;
        RECT 90.750 0.100 90.920 0.790 ;
        RECT 91.290 -0.070 91.460 0.800 ;
        RECT 91.730 0.760 92.150 1.040 ;
        RECT 93.370 0.930 93.540 1.260 ;
        RECT 92.670 0.760 94.090 0.930 ;
        RECT 91.730 0.320 93.310 0.490 ;
        RECT 88.560 -0.450 88.730 -0.120 ;
        RECT 89.970 -0.240 91.550 -0.070 ;
        RECT 87.030 -0.720 87.450 -0.510 ;
        RECT 87.920 -0.720 88.340 -0.510 ;
        RECT 89.150 -0.680 90.610 -0.510 ;
        RECT 87.100 -0.780 87.360 -0.720 ;
        RECT 88.010 -0.780 88.270 -0.720 ;
        RECT 89.610 -0.740 89.900 -0.680 ;
        RECT 91.130 -0.850 91.550 -0.510 ;
        RECT 91.810 -0.550 91.980 0.320 ;
        RECT 92.360 -0.550 92.530 0.140 ;
        RECT 94.310 -0.450 94.480 -0.120 ;
        RECT 92.780 -0.720 93.200 -0.510 ;
        RECT 93.670 -0.720 94.090 -0.510 ;
        RECT 92.850 -0.780 93.110 -0.720 ;
        RECT 93.760 -0.780 94.020 -0.720 ;
        RECT 2.990 -1.440 3.250 -1.350 ;
        RECT 3.900 -1.440 4.160 -1.350 ;
        RECT 2.900 -1.650 3.320 -1.440 ;
        RECT 3.830 -1.650 4.250 -1.440 ;
        RECT 2.520 -2.040 2.690 -1.710 ;
        RECT 4.500 -2.310 4.670 -1.620 ;
        RECT 5.040 -2.480 5.210 -1.610 ;
        RECT 5.480 -1.650 5.900 -1.370 ;
        RECT 7.120 -1.480 7.290 -1.150 ;
        RECT 8.740 -1.440 9.000 -1.350 ;
        RECT 9.650 -1.440 9.910 -1.350 ;
        RECT 6.420 -1.650 7.840 -1.480 ;
        RECT 8.650 -1.650 9.070 -1.440 ;
        RECT 9.580 -1.650 10.000 -1.440 ;
        RECT 5.480 -2.090 7.060 -1.920 ;
        RECT 8.270 -2.040 8.440 -1.710 ;
        RECT 3.720 -2.650 5.300 -2.480 ;
        RECT 2.900 -3.090 4.360 -2.920 ;
        RECT 3.360 -3.150 3.650 -3.090 ;
        RECT 4.880 -3.260 5.300 -2.920 ;
        RECT 5.560 -2.960 5.730 -2.090 ;
        RECT 6.110 -2.960 6.280 -2.270 ;
        RECT 10.250 -2.310 10.420 -1.620 ;
        RECT 10.790 -2.480 10.960 -1.610 ;
        RECT 11.230 -1.650 11.650 -1.370 ;
        RECT 12.870 -1.480 13.040 -1.150 ;
        RECT 14.490 -1.440 14.750 -1.350 ;
        RECT 15.400 -1.440 15.660 -1.350 ;
        RECT 12.170 -1.650 13.590 -1.480 ;
        RECT 14.400 -1.650 14.820 -1.440 ;
        RECT 15.330 -1.650 15.750 -1.440 ;
        RECT 11.230 -2.090 12.810 -1.920 ;
        RECT 14.020 -2.040 14.190 -1.710 ;
        RECT 8.060 -2.860 8.230 -2.530 ;
        RECT 9.470 -2.650 11.050 -2.480 ;
        RECT 6.530 -3.130 6.950 -2.920 ;
        RECT 7.420 -3.130 7.840 -2.920 ;
        RECT 8.650 -3.090 10.110 -2.920 ;
        RECT 6.600 -3.190 6.860 -3.130 ;
        RECT 7.510 -3.190 7.770 -3.130 ;
        RECT 9.110 -3.150 9.400 -3.090 ;
        RECT 10.630 -3.260 11.050 -2.920 ;
        RECT 11.310 -2.960 11.480 -2.090 ;
        RECT 11.860 -2.960 12.030 -2.270 ;
        RECT 16.000 -2.310 16.170 -1.620 ;
        RECT 16.540 -2.480 16.710 -1.610 ;
        RECT 16.980 -1.650 17.400 -1.370 ;
        RECT 18.620 -1.480 18.790 -1.150 ;
        RECT 20.240 -1.440 20.500 -1.350 ;
        RECT 21.150 -1.440 21.410 -1.350 ;
        RECT 17.920 -1.650 19.340 -1.480 ;
        RECT 20.150 -1.650 20.570 -1.440 ;
        RECT 21.080 -1.650 21.500 -1.440 ;
        RECT 16.980 -2.090 18.560 -1.920 ;
        RECT 19.770 -2.040 19.940 -1.710 ;
        RECT 13.810 -2.860 13.980 -2.530 ;
        RECT 15.220 -2.650 16.800 -2.480 ;
        RECT 12.280 -3.130 12.700 -2.920 ;
        RECT 13.170 -3.130 13.590 -2.920 ;
        RECT 14.400 -3.090 15.860 -2.920 ;
        RECT 12.350 -3.190 12.610 -3.130 ;
        RECT 13.260 -3.190 13.520 -3.130 ;
        RECT 14.860 -3.150 15.150 -3.090 ;
        RECT 16.380 -3.260 16.800 -2.920 ;
        RECT 17.060 -2.960 17.230 -2.090 ;
        RECT 17.610 -2.960 17.780 -2.270 ;
        RECT 21.750 -2.310 21.920 -1.620 ;
        RECT 22.290 -2.480 22.460 -1.610 ;
        RECT 22.730 -1.650 23.150 -1.370 ;
        RECT 24.370 -1.480 24.540 -1.150 ;
        RECT 25.990 -1.440 26.250 -1.350 ;
        RECT 26.900 -1.440 27.160 -1.350 ;
        RECT 23.670 -1.650 25.090 -1.480 ;
        RECT 25.900 -1.650 26.320 -1.440 ;
        RECT 26.830 -1.650 27.250 -1.440 ;
        RECT 22.730 -2.090 24.310 -1.920 ;
        RECT 25.520 -2.040 25.690 -1.710 ;
        RECT 19.560 -2.860 19.730 -2.530 ;
        RECT 20.970 -2.650 22.550 -2.480 ;
        RECT 18.030 -3.130 18.450 -2.920 ;
        RECT 18.920 -3.130 19.340 -2.920 ;
        RECT 20.150 -3.090 21.610 -2.920 ;
        RECT 18.100 -3.190 18.360 -3.130 ;
        RECT 19.010 -3.190 19.270 -3.130 ;
        RECT 20.610 -3.150 20.900 -3.090 ;
        RECT 22.130 -3.260 22.550 -2.920 ;
        RECT 22.810 -2.960 22.980 -2.090 ;
        RECT 23.360 -2.960 23.530 -2.270 ;
        RECT 27.500 -2.310 27.670 -1.620 ;
        RECT 28.040 -2.480 28.210 -1.610 ;
        RECT 28.480 -1.650 28.900 -1.370 ;
        RECT 30.120 -1.480 30.290 -1.150 ;
        RECT 31.740 -1.440 32.000 -1.350 ;
        RECT 32.650 -1.440 32.910 -1.350 ;
        RECT 29.420 -1.650 30.840 -1.480 ;
        RECT 31.650 -1.650 32.070 -1.440 ;
        RECT 32.580 -1.650 33.000 -1.440 ;
        RECT 28.480 -2.090 30.060 -1.920 ;
        RECT 31.270 -2.040 31.440 -1.710 ;
        RECT 25.310 -2.860 25.480 -2.530 ;
        RECT 26.720 -2.650 28.300 -2.480 ;
        RECT 23.780 -3.130 24.200 -2.920 ;
        RECT 24.670 -3.130 25.090 -2.920 ;
        RECT 25.900 -3.090 27.360 -2.920 ;
        RECT 23.850 -3.190 24.110 -3.130 ;
        RECT 24.760 -3.190 25.020 -3.130 ;
        RECT 26.360 -3.150 26.650 -3.090 ;
        RECT 27.880 -3.260 28.300 -2.920 ;
        RECT 28.560 -2.960 28.730 -2.090 ;
        RECT 29.110 -2.960 29.280 -2.270 ;
        RECT 33.250 -2.310 33.420 -1.620 ;
        RECT 33.790 -2.480 33.960 -1.610 ;
        RECT 34.230 -1.650 34.650 -1.370 ;
        RECT 35.870 -1.480 36.040 -1.150 ;
        RECT 37.490 -1.440 37.750 -1.350 ;
        RECT 38.400 -1.440 38.660 -1.350 ;
        RECT 35.170 -1.650 36.590 -1.480 ;
        RECT 37.400 -1.650 37.820 -1.440 ;
        RECT 38.330 -1.650 38.750 -1.440 ;
        RECT 34.230 -2.090 35.810 -1.920 ;
        RECT 37.020 -2.040 37.190 -1.710 ;
        RECT 31.060 -2.860 31.230 -2.530 ;
        RECT 32.470 -2.650 34.050 -2.480 ;
        RECT 29.530 -3.130 29.950 -2.920 ;
        RECT 30.420 -3.130 30.840 -2.920 ;
        RECT 31.650 -3.090 33.110 -2.920 ;
        RECT 29.600 -3.190 29.860 -3.130 ;
        RECT 30.510 -3.190 30.770 -3.130 ;
        RECT 32.110 -3.150 32.400 -3.090 ;
        RECT 33.630 -3.260 34.050 -2.920 ;
        RECT 34.310 -2.960 34.480 -2.090 ;
        RECT 34.860 -2.960 35.030 -2.270 ;
        RECT 39.000 -2.310 39.170 -1.620 ;
        RECT 39.540 -2.480 39.710 -1.610 ;
        RECT 39.980 -1.650 40.400 -1.370 ;
        RECT 41.620 -1.480 41.790 -1.150 ;
        RECT 43.240 -1.440 43.500 -1.350 ;
        RECT 44.150 -1.440 44.410 -1.350 ;
        RECT 40.920 -1.650 42.340 -1.480 ;
        RECT 43.150 -1.650 43.570 -1.440 ;
        RECT 44.080 -1.650 44.500 -1.440 ;
        RECT 39.980 -2.090 41.560 -1.920 ;
        RECT 42.770 -2.040 42.940 -1.710 ;
        RECT 36.810 -2.860 36.980 -2.530 ;
        RECT 38.220 -2.650 39.800 -2.480 ;
        RECT 35.280 -3.130 35.700 -2.920 ;
        RECT 36.170 -3.130 36.590 -2.920 ;
        RECT 37.400 -3.090 38.860 -2.920 ;
        RECT 35.350 -3.190 35.610 -3.130 ;
        RECT 36.260 -3.190 36.520 -3.130 ;
        RECT 37.860 -3.150 38.150 -3.090 ;
        RECT 39.380 -3.260 39.800 -2.920 ;
        RECT 40.060 -2.960 40.230 -2.090 ;
        RECT 40.610 -2.960 40.780 -2.270 ;
        RECT 44.750 -2.310 44.920 -1.620 ;
        RECT 45.290 -2.480 45.460 -1.610 ;
        RECT 45.730 -1.650 46.150 -1.370 ;
        RECT 47.370 -1.480 47.540 -1.150 ;
        RECT 48.990 -1.440 49.250 -1.350 ;
        RECT 49.900 -1.440 50.160 -1.350 ;
        RECT 46.670 -1.650 48.090 -1.480 ;
        RECT 48.900 -1.650 49.320 -1.440 ;
        RECT 49.830 -1.650 50.250 -1.440 ;
        RECT 45.730 -2.090 47.310 -1.920 ;
        RECT 48.520 -2.040 48.690 -1.710 ;
        RECT 42.560 -2.860 42.730 -2.530 ;
        RECT 43.970 -2.650 45.550 -2.480 ;
        RECT 41.030 -3.130 41.450 -2.920 ;
        RECT 41.920 -3.130 42.340 -2.920 ;
        RECT 43.150 -3.090 44.610 -2.920 ;
        RECT 41.100 -3.190 41.360 -3.130 ;
        RECT 42.010 -3.190 42.270 -3.130 ;
        RECT 43.610 -3.150 43.900 -3.090 ;
        RECT 45.130 -3.260 45.550 -2.920 ;
        RECT 45.810 -2.960 45.980 -2.090 ;
        RECT 46.360 -2.960 46.530 -2.270 ;
        RECT 50.500 -2.310 50.670 -1.620 ;
        RECT 51.040 -2.480 51.210 -1.610 ;
        RECT 51.480 -1.650 51.900 -1.370 ;
        RECT 53.120 -1.480 53.290 -1.150 ;
        RECT 54.740 -1.440 55.000 -1.350 ;
        RECT 55.650 -1.440 55.910 -1.350 ;
        RECT 52.420 -1.650 53.840 -1.480 ;
        RECT 54.650 -1.650 55.070 -1.440 ;
        RECT 55.580 -1.650 56.000 -1.440 ;
        RECT 51.480 -2.090 53.060 -1.920 ;
        RECT 54.270 -2.040 54.440 -1.710 ;
        RECT 48.310 -2.860 48.480 -2.530 ;
        RECT 49.720 -2.650 51.300 -2.480 ;
        RECT 46.780 -3.130 47.200 -2.920 ;
        RECT 47.670 -3.130 48.090 -2.920 ;
        RECT 48.900 -3.090 50.360 -2.920 ;
        RECT 46.850 -3.190 47.110 -3.130 ;
        RECT 47.760 -3.190 48.020 -3.130 ;
        RECT 49.360 -3.150 49.650 -3.090 ;
        RECT 50.880 -3.260 51.300 -2.920 ;
        RECT 51.560 -2.960 51.730 -2.090 ;
        RECT 52.110 -2.960 52.280 -2.270 ;
        RECT 56.250 -2.310 56.420 -1.620 ;
        RECT 56.790 -2.480 56.960 -1.610 ;
        RECT 57.230 -1.650 57.650 -1.370 ;
        RECT 58.870 -1.480 59.040 -1.150 ;
        RECT 60.490 -1.440 60.750 -1.350 ;
        RECT 61.400 -1.440 61.660 -1.350 ;
        RECT 58.170 -1.650 59.590 -1.480 ;
        RECT 60.400 -1.650 60.820 -1.440 ;
        RECT 61.330 -1.650 61.750 -1.440 ;
        RECT 57.230 -2.090 58.810 -1.920 ;
        RECT 60.020 -2.040 60.190 -1.710 ;
        RECT 54.060 -2.860 54.230 -2.530 ;
        RECT 55.470 -2.650 57.050 -2.480 ;
        RECT 52.530 -3.130 52.950 -2.920 ;
        RECT 53.420 -3.130 53.840 -2.920 ;
        RECT 54.650 -3.090 56.110 -2.920 ;
        RECT 52.600 -3.190 52.860 -3.130 ;
        RECT 53.510 -3.190 53.770 -3.130 ;
        RECT 55.110 -3.150 55.400 -3.090 ;
        RECT 56.630 -3.260 57.050 -2.920 ;
        RECT 57.310 -2.960 57.480 -2.090 ;
        RECT 57.860 -2.960 58.030 -2.270 ;
        RECT 62.000 -2.310 62.170 -1.620 ;
        RECT 62.540 -2.480 62.710 -1.610 ;
        RECT 62.980 -1.650 63.400 -1.370 ;
        RECT 64.620 -1.480 64.790 -1.150 ;
        RECT 66.240 -1.440 66.500 -1.350 ;
        RECT 67.150 -1.440 67.410 -1.350 ;
        RECT 63.920 -1.650 65.340 -1.480 ;
        RECT 66.150 -1.650 66.570 -1.440 ;
        RECT 67.080 -1.650 67.500 -1.440 ;
        RECT 62.980 -2.090 64.560 -1.920 ;
        RECT 65.770 -2.040 65.940 -1.710 ;
        RECT 59.810 -2.860 59.980 -2.530 ;
        RECT 61.220 -2.650 62.800 -2.480 ;
        RECT 58.280 -3.130 58.700 -2.920 ;
        RECT 59.170 -3.130 59.590 -2.920 ;
        RECT 60.400 -3.090 61.860 -2.920 ;
        RECT 58.350 -3.190 58.610 -3.130 ;
        RECT 59.260 -3.190 59.520 -3.130 ;
        RECT 60.860 -3.150 61.150 -3.090 ;
        RECT 62.380 -3.260 62.800 -2.920 ;
        RECT 63.060 -2.960 63.230 -2.090 ;
        RECT 63.610 -2.960 63.780 -2.270 ;
        RECT 67.750 -2.310 67.920 -1.620 ;
        RECT 68.290 -2.480 68.460 -1.610 ;
        RECT 68.730 -1.650 69.150 -1.370 ;
        RECT 70.370 -1.480 70.540 -1.150 ;
        RECT 71.990 -1.440 72.250 -1.350 ;
        RECT 72.900 -1.440 73.160 -1.350 ;
        RECT 69.670 -1.650 71.090 -1.480 ;
        RECT 71.900 -1.650 72.320 -1.440 ;
        RECT 72.830 -1.650 73.250 -1.440 ;
        RECT 68.730 -2.090 70.310 -1.920 ;
        RECT 71.520 -2.040 71.690 -1.710 ;
        RECT 65.560 -2.860 65.730 -2.530 ;
        RECT 66.970 -2.650 68.550 -2.480 ;
        RECT 64.030 -3.130 64.450 -2.920 ;
        RECT 64.920 -3.130 65.340 -2.920 ;
        RECT 66.150 -3.090 67.610 -2.920 ;
        RECT 64.100 -3.190 64.360 -3.130 ;
        RECT 65.010 -3.190 65.270 -3.130 ;
        RECT 66.610 -3.150 66.900 -3.090 ;
        RECT 68.130 -3.260 68.550 -2.920 ;
        RECT 68.810 -2.960 68.980 -2.090 ;
        RECT 69.360 -2.960 69.530 -2.270 ;
        RECT 73.500 -2.310 73.670 -1.620 ;
        RECT 74.040 -2.480 74.210 -1.610 ;
        RECT 74.480 -1.650 74.900 -1.370 ;
        RECT 76.120 -1.480 76.290 -1.150 ;
        RECT 77.740 -1.440 78.000 -1.350 ;
        RECT 78.650 -1.440 78.910 -1.350 ;
        RECT 75.420 -1.650 76.840 -1.480 ;
        RECT 77.650 -1.650 78.070 -1.440 ;
        RECT 78.580 -1.650 79.000 -1.440 ;
        RECT 74.480 -2.090 76.060 -1.920 ;
        RECT 77.270 -2.040 77.440 -1.710 ;
        RECT 71.310 -2.860 71.480 -2.530 ;
        RECT 72.720 -2.650 74.300 -2.480 ;
        RECT 69.780 -3.130 70.200 -2.920 ;
        RECT 70.670 -3.130 71.090 -2.920 ;
        RECT 71.900 -3.090 73.360 -2.920 ;
        RECT 69.850 -3.190 70.110 -3.130 ;
        RECT 70.760 -3.190 71.020 -3.130 ;
        RECT 72.360 -3.150 72.650 -3.090 ;
        RECT 73.880 -3.260 74.300 -2.920 ;
        RECT 74.560 -2.960 74.730 -2.090 ;
        RECT 75.110 -2.960 75.280 -2.270 ;
        RECT 79.250 -2.310 79.420 -1.620 ;
        RECT 79.790 -2.480 79.960 -1.610 ;
        RECT 80.230 -1.650 80.650 -1.370 ;
        RECT 81.870 -1.480 82.040 -1.150 ;
        RECT 83.490 -1.440 83.750 -1.350 ;
        RECT 84.400 -1.440 84.660 -1.350 ;
        RECT 81.170 -1.650 82.590 -1.480 ;
        RECT 83.400 -1.650 83.820 -1.440 ;
        RECT 84.330 -1.650 84.750 -1.440 ;
        RECT 80.230 -2.090 81.810 -1.920 ;
        RECT 83.020 -2.040 83.190 -1.710 ;
        RECT 77.060 -2.860 77.230 -2.530 ;
        RECT 78.470 -2.650 80.050 -2.480 ;
        RECT 75.530 -3.130 75.950 -2.920 ;
        RECT 76.420 -3.130 76.840 -2.920 ;
        RECT 77.650 -3.090 79.110 -2.920 ;
        RECT 75.600 -3.190 75.860 -3.130 ;
        RECT 76.510 -3.190 76.770 -3.130 ;
        RECT 78.110 -3.150 78.400 -3.090 ;
        RECT 79.630 -3.260 80.050 -2.920 ;
        RECT 80.310 -2.960 80.480 -2.090 ;
        RECT 80.860 -2.960 81.030 -2.270 ;
        RECT 85.000 -2.310 85.170 -1.620 ;
        RECT 85.540 -2.480 85.710 -1.610 ;
        RECT 85.980 -1.650 86.400 -1.370 ;
        RECT 87.620 -1.480 87.790 -1.150 ;
        RECT 89.240 -1.440 89.500 -1.350 ;
        RECT 90.150 -1.440 90.410 -1.350 ;
        RECT 86.920 -1.650 88.340 -1.480 ;
        RECT 89.150 -1.650 89.570 -1.440 ;
        RECT 90.080 -1.650 90.500 -1.440 ;
        RECT 85.980 -2.090 87.560 -1.920 ;
        RECT 88.770 -2.040 88.940 -1.710 ;
        RECT 82.810 -2.860 82.980 -2.530 ;
        RECT 84.220 -2.650 85.800 -2.480 ;
        RECT 81.280 -3.130 81.700 -2.920 ;
        RECT 82.170 -3.130 82.590 -2.920 ;
        RECT 83.400 -3.090 84.860 -2.920 ;
        RECT 81.350 -3.190 81.610 -3.130 ;
        RECT 82.260 -3.190 82.520 -3.130 ;
        RECT 83.860 -3.150 84.150 -3.090 ;
        RECT 85.380 -3.260 85.800 -2.920 ;
        RECT 86.060 -2.960 86.230 -2.090 ;
        RECT 86.610 -2.960 86.780 -2.270 ;
        RECT 90.750 -2.310 90.920 -1.620 ;
        RECT 91.290 -2.480 91.460 -1.610 ;
        RECT 91.730 -1.650 92.150 -1.370 ;
        RECT 93.370 -1.480 93.540 -1.150 ;
        RECT 92.670 -1.650 94.090 -1.480 ;
        RECT 91.730 -2.090 93.310 -1.920 ;
        RECT 88.560 -2.860 88.730 -2.530 ;
        RECT 89.970 -2.650 91.550 -2.480 ;
        RECT 87.030 -3.130 87.450 -2.920 ;
        RECT 87.920 -3.130 88.340 -2.920 ;
        RECT 89.150 -3.090 90.610 -2.920 ;
        RECT 87.100 -3.190 87.360 -3.130 ;
        RECT 88.010 -3.190 88.270 -3.130 ;
        RECT 89.610 -3.150 89.900 -3.090 ;
        RECT 91.130 -3.260 91.550 -2.920 ;
        RECT 91.810 -2.960 91.980 -2.090 ;
        RECT 92.360 -2.960 92.530 -2.270 ;
        RECT 94.310 -2.860 94.480 -2.530 ;
        RECT 92.780 -3.130 93.200 -2.920 ;
        RECT 93.670 -3.130 94.090 -2.920 ;
        RECT 92.850 -3.190 93.110 -3.130 ;
        RECT 93.760 -3.190 94.020 -3.130 ;
        RECT 2.990 -3.850 3.250 -3.760 ;
        RECT 3.900 -3.850 4.160 -3.760 ;
        RECT 2.900 -4.060 3.320 -3.850 ;
        RECT 3.830 -4.060 4.250 -3.850 ;
        RECT 2.520 -4.450 2.690 -4.120 ;
        RECT 4.500 -4.720 4.670 -4.030 ;
        RECT 5.040 -4.890 5.210 -4.020 ;
        RECT 5.480 -4.060 5.900 -3.780 ;
        RECT 7.120 -3.890 7.290 -3.560 ;
        RECT 8.740 -3.850 9.000 -3.760 ;
        RECT 9.650 -3.850 9.910 -3.760 ;
        RECT 6.420 -4.060 7.840 -3.890 ;
        RECT 8.650 -4.060 9.070 -3.850 ;
        RECT 9.580 -4.060 10.000 -3.850 ;
        RECT 5.480 -4.500 7.060 -4.330 ;
        RECT 8.270 -4.450 8.440 -4.120 ;
        RECT 3.720 -5.060 5.300 -4.890 ;
        RECT 2.900 -5.500 4.360 -5.330 ;
        RECT 3.020 -6.380 3.190 -5.500 ;
        RECT 3.360 -5.560 3.650 -5.500 ;
        RECT 4.880 -5.670 5.300 -5.330 ;
        RECT 5.560 -5.370 5.730 -4.500 ;
        RECT 6.110 -5.370 6.280 -4.680 ;
        RECT 10.250 -4.720 10.420 -4.030 ;
        RECT 10.790 -4.890 10.960 -4.020 ;
        RECT 11.230 -4.060 11.650 -3.780 ;
        RECT 12.870 -3.890 13.040 -3.560 ;
        RECT 14.490 -3.850 14.750 -3.760 ;
        RECT 15.400 -3.850 15.660 -3.760 ;
        RECT 12.170 -4.060 13.590 -3.890 ;
        RECT 14.400 -4.060 14.820 -3.850 ;
        RECT 15.330 -4.060 15.750 -3.850 ;
        RECT 11.230 -4.500 12.810 -4.330 ;
        RECT 14.020 -4.450 14.190 -4.120 ;
        RECT 8.060 -5.270 8.230 -4.940 ;
        RECT 9.470 -5.060 11.050 -4.890 ;
        RECT 6.530 -5.540 6.950 -5.330 ;
        RECT 7.420 -5.540 7.840 -5.330 ;
        RECT 8.650 -5.500 10.110 -5.330 ;
        RECT 6.600 -5.600 6.860 -5.540 ;
        RECT 7.510 -5.600 7.770 -5.540 ;
        RECT 5.010 -6.380 5.180 -5.670 ;
        RECT 2.990 -6.850 3.250 -6.760 ;
        RECT 3.900 -6.850 4.160 -6.760 ;
        RECT 2.900 -7.060 3.320 -6.850 ;
        RECT 3.830 -7.060 4.250 -6.850 ;
        RECT 2.520 -7.450 2.690 -7.120 ;
        RECT 4.500 -7.720 4.670 -7.030 ;
        RECT 5.040 -7.890 5.210 -7.020 ;
        RECT 5.480 -7.060 5.900 -6.780 ;
        RECT 7.120 -6.890 7.290 -6.290 ;
        RECT 8.770 -6.380 8.940 -5.500 ;
        RECT 9.110 -5.560 9.400 -5.500 ;
        RECT 10.630 -5.670 11.050 -5.330 ;
        RECT 11.310 -5.370 11.480 -4.500 ;
        RECT 11.860 -5.370 12.030 -4.680 ;
        RECT 16.000 -4.720 16.170 -4.030 ;
        RECT 16.540 -4.890 16.710 -4.020 ;
        RECT 16.980 -4.060 17.400 -3.780 ;
        RECT 18.620 -3.890 18.790 -3.560 ;
        RECT 20.240 -3.850 20.500 -3.760 ;
        RECT 21.150 -3.850 21.410 -3.760 ;
        RECT 17.920 -4.060 19.340 -3.890 ;
        RECT 20.150 -4.060 20.570 -3.850 ;
        RECT 21.080 -4.060 21.500 -3.850 ;
        RECT 16.980 -4.500 18.560 -4.330 ;
        RECT 19.770 -4.450 19.940 -4.120 ;
        RECT 13.810 -5.270 13.980 -4.940 ;
        RECT 15.220 -5.060 16.800 -4.890 ;
        RECT 12.280 -5.540 12.700 -5.330 ;
        RECT 13.170 -5.540 13.590 -5.330 ;
        RECT 14.400 -5.500 15.860 -5.330 ;
        RECT 12.350 -5.600 12.610 -5.540 ;
        RECT 13.260 -5.600 13.520 -5.540 ;
        RECT 10.770 -6.380 10.940 -5.670 ;
        RECT 8.740 -6.850 9.000 -6.760 ;
        RECT 9.650 -6.850 9.910 -6.760 ;
        RECT 6.420 -7.060 7.840 -6.890 ;
        RECT 8.650 -7.060 9.070 -6.850 ;
        RECT 9.580 -7.060 10.000 -6.850 ;
        RECT 5.480 -7.500 7.060 -7.330 ;
        RECT 8.270 -7.450 8.440 -7.120 ;
        RECT 3.720 -8.060 5.300 -7.890 ;
        RECT 2.900 -8.500 4.360 -8.330 ;
        RECT 3.360 -8.560 3.650 -8.500 ;
        RECT 4.880 -8.670 5.300 -8.330 ;
        RECT 5.560 -8.370 5.730 -7.500 ;
        RECT 6.110 -8.370 6.280 -7.680 ;
        RECT 10.250 -7.720 10.420 -7.030 ;
        RECT 10.790 -7.890 10.960 -7.020 ;
        RECT 11.230 -7.060 11.650 -6.780 ;
        RECT 12.870 -6.890 13.040 -6.290 ;
        RECT 14.520 -6.380 14.690 -5.500 ;
        RECT 14.860 -5.560 15.150 -5.500 ;
        RECT 16.380 -5.670 16.800 -5.330 ;
        RECT 17.060 -5.370 17.230 -4.500 ;
        RECT 17.610 -5.370 17.780 -4.680 ;
        RECT 21.750 -4.720 21.920 -4.030 ;
        RECT 22.290 -4.890 22.460 -4.020 ;
        RECT 22.730 -4.060 23.150 -3.780 ;
        RECT 24.370 -3.890 24.540 -3.560 ;
        RECT 25.990 -3.850 26.250 -3.760 ;
        RECT 26.900 -3.850 27.160 -3.760 ;
        RECT 23.670 -4.060 25.090 -3.890 ;
        RECT 25.900 -4.060 26.320 -3.850 ;
        RECT 26.830 -4.060 27.250 -3.850 ;
        RECT 22.730 -4.500 24.310 -4.330 ;
        RECT 25.520 -4.450 25.690 -4.120 ;
        RECT 19.560 -5.270 19.730 -4.940 ;
        RECT 20.970 -5.060 22.550 -4.890 ;
        RECT 18.030 -5.540 18.450 -5.330 ;
        RECT 18.920 -5.540 19.340 -5.330 ;
        RECT 20.150 -5.500 21.610 -5.330 ;
        RECT 18.100 -5.600 18.360 -5.540 ;
        RECT 19.010 -5.600 19.270 -5.540 ;
        RECT 16.520 -6.380 16.690 -5.670 ;
        RECT 14.490 -6.850 14.750 -6.760 ;
        RECT 15.400 -6.850 15.660 -6.760 ;
        RECT 12.170 -7.060 13.590 -6.890 ;
        RECT 14.400 -7.060 14.820 -6.850 ;
        RECT 15.330 -7.060 15.750 -6.850 ;
        RECT 11.230 -7.500 12.810 -7.330 ;
        RECT 14.020 -7.450 14.190 -7.120 ;
        RECT 8.060 -8.270 8.230 -7.940 ;
        RECT 9.470 -8.060 11.050 -7.890 ;
        RECT 6.530 -8.540 6.950 -8.330 ;
        RECT 7.420 -8.540 7.840 -8.330 ;
        RECT 8.650 -8.500 10.110 -8.330 ;
        RECT 6.600 -8.600 6.860 -8.540 ;
        RECT 7.510 -8.600 7.770 -8.540 ;
        RECT 9.110 -8.560 9.400 -8.500 ;
        RECT 10.630 -8.670 11.050 -8.330 ;
        RECT 11.310 -8.370 11.480 -7.500 ;
        RECT 11.860 -8.370 12.030 -7.680 ;
        RECT 16.000 -7.720 16.170 -7.030 ;
        RECT 16.540 -7.890 16.710 -7.020 ;
        RECT 16.980 -7.060 17.400 -6.780 ;
        RECT 18.620 -6.890 18.790 -6.290 ;
        RECT 20.270 -6.380 20.440 -5.500 ;
        RECT 20.610 -5.560 20.900 -5.500 ;
        RECT 22.130 -5.670 22.550 -5.330 ;
        RECT 22.810 -5.370 22.980 -4.500 ;
        RECT 23.360 -5.370 23.530 -4.680 ;
        RECT 27.500 -4.720 27.670 -4.030 ;
        RECT 28.040 -4.890 28.210 -4.020 ;
        RECT 28.480 -4.060 28.900 -3.780 ;
        RECT 30.120 -3.890 30.290 -3.560 ;
        RECT 31.740 -3.850 32.000 -3.760 ;
        RECT 32.650 -3.850 32.910 -3.760 ;
        RECT 29.420 -4.060 30.840 -3.890 ;
        RECT 31.650 -4.060 32.070 -3.850 ;
        RECT 32.580 -4.060 33.000 -3.850 ;
        RECT 28.480 -4.500 30.060 -4.330 ;
        RECT 31.270 -4.450 31.440 -4.120 ;
        RECT 25.310 -5.270 25.480 -4.940 ;
        RECT 26.720 -5.060 28.300 -4.890 ;
        RECT 23.780 -5.540 24.200 -5.330 ;
        RECT 24.670 -5.540 25.090 -5.330 ;
        RECT 25.900 -5.500 27.360 -5.330 ;
        RECT 23.850 -5.600 24.110 -5.540 ;
        RECT 24.760 -5.600 25.020 -5.540 ;
        RECT 22.270 -6.380 22.440 -5.670 ;
        RECT 20.240 -6.850 20.500 -6.760 ;
        RECT 21.150 -6.850 21.410 -6.760 ;
        RECT 17.920 -7.060 19.340 -6.890 ;
        RECT 20.150 -7.060 20.570 -6.850 ;
        RECT 21.080 -7.060 21.500 -6.850 ;
        RECT 16.980 -7.500 18.560 -7.330 ;
        RECT 19.770 -7.450 19.940 -7.120 ;
        RECT 13.810 -8.270 13.980 -7.940 ;
        RECT 15.220 -8.060 16.800 -7.890 ;
        RECT 12.280 -8.540 12.700 -8.330 ;
        RECT 13.170 -8.540 13.590 -8.330 ;
        RECT 14.400 -8.500 15.860 -8.330 ;
        RECT 12.350 -8.600 12.610 -8.540 ;
        RECT 13.260 -8.600 13.520 -8.540 ;
        RECT 14.860 -8.560 15.150 -8.500 ;
        RECT 16.380 -8.670 16.800 -8.330 ;
        RECT 17.060 -8.370 17.230 -7.500 ;
        RECT 17.610 -8.370 17.780 -7.680 ;
        RECT 21.750 -7.720 21.920 -7.030 ;
        RECT 22.290 -7.890 22.460 -7.020 ;
        RECT 22.730 -7.060 23.150 -6.780 ;
        RECT 24.370 -6.890 24.540 -6.290 ;
        RECT 26.020 -6.380 26.190 -5.500 ;
        RECT 26.360 -5.560 26.650 -5.500 ;
        RECT 27.880 -5.670 28.300 -5.330 ;
        RECT 28.560 -5.370 28.730 -4.500 ;
        RECT 29.110 -5.370 29.280 -4.680 ;
        RECT 33.250 -4.720 33.420 -4.030 ;
        RECT 33.790 -4.890 33.960 -4.020 ;
        RECT 34.230 -4.060 34.650 -3.780 ;
        RECT 35.870 -3.890 36.040 -3.560 ;
        RECT 37.490 -3.850 37.750 -3.760 ;
        RECT 38.400 -3.850 38.660 -3.760 ;
        RECT 35.170 -4.060 36.590 -3.890 ;
        RECT 37.400 -4.060 37.820 -3.850 ;
        RECT 38.330 -4.060 38.750 -3.850 ;
        RECT 34.230 -4.500 35.810 -4.330 ;
        RECT 37.020 -4.450 37.190 -4.120 ;
        RECT 31.060 -5.270 31.230 -4.940 ;
        RECT 32.470 -5.060 34.050 -4.890 ;
        RECT 29.530 -5.540 29.950 -5.330 ;
        RECT 30.420 -5.540 30.840 -5.330 ;
        RECT 31.650 -5.500 33.110 -5.330 ;
        RECT 29.600 -5.600 29.860 -5.540 ;
        RECT 30.510 -5.600 30.770 -5.540 ;
        RECT 28.020 -6.380 28.190 -5.670 ;
        RECT 25.990 -6.850 26.250 -6.760 ;
        RECT 26.900 -6.850 27.160 -6.760 ;
        RECT 23.670 -7.060 25.090 -6.890 ;
        RECT 25.900 -7.060 26.320 -6.850 ;
        RECT 26.830 -7.060 27.250 -6.850 ;
        RECT 22.730 -7.500 24.310 -7.330 ;
        RECT 25.520 -7.450 25.690 -7.120 ;
        RECT 19.560 -8.270 19.730 -7.940 ;
        RECT 20.970 -8.060 22.550 -7.890 ;
        RECT 18.030 -8.540 18.450 -8.330 ;
        RECT 18.920 -8.540 19.340 -8.330 ;
        RECT 20.150 -8.500 21.610 -8.330 ;
        RECT 18.100 -8.600 18.360 -8.540 ;
        RECT 19.010 -8.600 19.270 -8.540 ;
        RECT 20.610 -8.560 20.900 -8.500 ;
        RECT 22.130 -8.670 22.550 -8.330 ;
        RECT 22.810 -8.370 22.980 -7.500 ;
        RECT 23.360 -8.370 23.530 -7.680 ;
        RECT 27.500 -7.720 27.670 -7.030 ;
        RECT 28.040 -7.890 28.210 -7.020 ;
        RECT 28.480 -7.060 28.900 -6.780 ;
        RECT 30.120 -6.890 30.290 -6.290 ;
        RECT 31.770 -6.380 31.940 -5.500 ;
        RECT 32.110 -5.560 32.400 -5.500 ;
        RECT 33.630 -5.670 34.050 -5.330 ;
        RECT 34.310 -5.370 34.480 -4.500 ;
        RECT 34.860 -5.370 35.030 -4.680 ;
        RECT 39.000 -4.720 39.170 -4.030 ;
        RECT 39.540 -4.890 39.710 -4.020 ;
        RECT 39.980 -4.060 40.400 -3.780 ;
        RECT 41.620 -3.890 41.790 -3.560 ;
        RECT 43.240 -3.850 43.500 -3.760 ;
        RECT 44.150 -3.850 44.410 -3.760 ;
        RECT 40.920 -4.060 42.340 -3.890 ;
        RECT 43.150 -4.060 43.570 -3.850 ;
        RECT 44.080 -4.060 44.500 -3.850 ;
        RECT 39.980 -4.500 41.560 -4.330 ;
        RECT 42.770 -4.450 42.940 -4.120 ;
        RECT 36.810 -5.270 36.980 -4.940 ;
        RECT 38.220 -5.060 39.800 -4.890 ;
        RECT 35.280 -5.540 35.700 -5.330 ;
        RECT 36.170 -5.540 36.590 -5.330 ;
        RECT 37.400 -5.500 38.860 -5.330 ;
        RECT 35.350 -5.600 35.610 -5.540 ;
        RECT 36.260 -5.600 36.520 -5.540 ;
        RECT 33.770 -6.380 33.940 -5.670 ;
        RECT 31.740 -6.850 32.000 -6.760 ;
        RECT 32.650 -6.850 32.910 -6.760 ;
        RECT 29.420 -7.060 30.840 -6.890 ;
        RECT 31.650 -7.060 32.070 -6.850 ;
        RECT 32.580 -7.060 33.000 -6.850 ;
        RECT 28.480 -7.500 30.060 -7.330 ;
        RECT 31.270 -7.450 31.440 -7.120 ;
        RECT 25.310 -8.270 25.480 -7.940 ;
        RECT 26.720 -8.060 28.300 -7.890 ;
        RECT 23.780 -8.540 24.200 -8.330 ;
        RECT 24.670 -8.540 25.090 -8.330 ;
        RECT 25.900 -8.500 27.360 -8.330 ;
        RECT 23.850 -8.600 24.110 -8.540 ;
        RECT 24.760 -8.600 25.020 -8.540 ;
        RECT 26.360 -8.560 26.650 -8.500 ;
        RECT 27.880 -8.670 28.300 -8.330 ;
        RECT 28.560 -8.370 28.730 -7.500 ;
        RECT 29.110 -8.370 29.280 -7.680 ;
        RECT 33.250 -7.720 33.420 -7.030 ;
        RECT 33.790 -7.890 33.960 -7.020 ;
        RECT 34.230 -7.060 34.650 -6.780 ;
        RECT 35.870 -6.890 36.040 -6.290 ;
        RECT 37.520 -6.380 37.690 -5.500 ;
        RECT 37.860 -5.560 38.150 -5.500 ;
        RECT 39.380 -5.670 39.800 -5.330 ;
        RECT 40.060 -5.370 40.230 -4.500 ;
        RECT 40.610 -5.370 40.780 -4.680 ;
        RECT 44.750 -4.720 44.920 -4.030 ;
        RECT 45.290 -4.890 45.460 -4.020 ;
        RECT 45.730 -4.060 46.150 -3.780 ;
        RECT 47.370 -3.890 47.540 -3.560 ;
        RECT 48.990 -3.850 49.250 -3.760 ;
        RECT 49.900 -3.850 50.160 -3.760 ;
        RECT 46.670 -4.060 48.090 -3.890 ;
        RECT 48.900 -4.060 49.320 -3.850 ;
        RECT 49.830 -4.060 50.250 -3.850 ;
        RECT 45.730 -4.500 47.310 -4.330 ;
        RECT 48.520 -4.450 48.690 -4.120 ;
        RECT 42.560 -5.270 42.730 -4.940 ;
        RECT 43.970 -5.060 45.550 -4.890 ;
        RECT 41.030 -5.540 41.450 -5.330 ;
        RECT 41.920 -5.540 42.340 -5.330 ;
        RECT 43.150 -5.500 44.610 -5.330 ;
        RECT 41.100 -5.600 41.360 -5.540 ;
        RECT 42.010 -5.600 42.270 -5.540 ;
        RECT 39.520 -6.380 39.690 -5.670 ;
        RECT 37.490 -6.850 37.750 -6.760 ;
        RECT 38.400 -6.850 38.660 -6.760 ;
        RECT 35.170 -7.060 36.590 -6.890 ;
        RECT 37.400 -7.060 37.820 -6.850 ;
        RECT 38.330 -7.060 38.750 -6.850 ;
        RECT 34.230 -7.500 35.810 -7.330 ;
        RECT 37.020 -7.450 37.190 -7.120 ;
        RECT 31.060 -8.270 31.230 -7.940 ;
        RECT 32.470 -8.060 34.050 -7.890 ;
        RECT 29.530 -8.540 29.950 -8.330 ;
        RECT 30.420 -8.540 30.840 -8.330 ;
        RECT 31.650 -8.500 33.110 -8.330 ;
        RECT 29.600 -8.600 29.860 -8.540 ;
        RECT 30.510 -8.600 30.770 -8.540 ;
        RECT 32.110 -8.560 32.400 -8.500 ;
        RECT 33.630 -8.670 34.050 -8.330 ;
        RECT 34.310 -8.370 34.480 -7.500 ;
        RECT 34.860 -8.370 35.030 -7.680 ;
        RECT 39.000 -7.720 39.170 -7.030 ;
        RECT 39.540 -7.890 39.710 -7.020 ;
        RECT 39.980 -7.060 40.400 -6.780 ;
        RECT 41.620 -6.890 41.790 -6.290 ;
        RECT 43.270 -6.380 43.440 -5.500 ;
        RECT 43.610 -5.560 43.900 -5.500 ;
        RECT 45.130 -5.670 45.550 -5.330 ;
        RECT 45.810 -5.370 45.980 -4.500 ;
        RECT 46.360 -5.370 46.530 -4.680 ;
        RECT 50.500 -4.720 50.670 -4.030 ;
        RECT 51.040 -4.890 51.210 -4.020 ;
        RECT 51.480 -4.060 51.900 -3.780 ;
        RECT 53.120 -3.890 53.290 -3.560 ;
        RECT 54.740 -3.850 55.000 -3.760 ;
        RECT 55.650 -3.850 55.910 -3.760 ;
        RECT 52.420 -4.060 53.840 -3.890 ;
        RECT 54.650 -4.060 55.070 -3.850 ;
        RECT 55.580 -4.060 56.000 -3.850 ;
        RECT 51.480 -4.500 53.060 -4.330 ;
        RECT 54.270 -4.450 54.440 -4.120 ;
        RECT 48.310 -5.270 48.480 -4.940 ;
        RECT 49.720 -5.060 51.300 -4.890 ;
        RECT 46.780 -5.540 47.200 -5.330 ;
        RECT 47.670 -5.540 48.090 -5.330 ;
        RECT 48.900 -5.500 50.360 -5.330 ;
        RECT 46.850 -5.600 47.110 -5.540 ;
        RECT 47.760 -5.600 48.020 -5.540 ;
        RECT 45.270 -6.380 45.440 -5.670 ;
        RECT 43.240 -6.850 43.500 -6.760 ;
        RECT 44.150 -6.850 44.410 -6.760 ;
        RECT 40.920 -7.060 42.340 -6.890 ;
        RECT 43.150 -7.060 43.570 -6.850 ;
        RECT 44.080 -7.060 44.500 -6.850 ;
        RECT 39.980 -7.500 41.560 -7.330 ;
        RECT 42.770 -7.450 42.940 -7.120 ;
        RECT 36.810 -8.270 36.980 -7.940 ;
        RECT 38.220 -8.060 39.800 -7.890 ;
        RECT 35.280 -8.540 35.700 -8.330 ;
        RECT 36.170 -8.540 36.590 -8.330 ;
        RECT 37.400 -8.500 38.860 -8.330 ;
        RECT 35.350 -8.600 35.610 -8.540 ;
        RECT 36.260 -8.600 36.520 -8.540 ;
        RECT 37.860 -8.560 38.150 -8.500 ;
        RECT 39.380 -8.670 39.800 -8.330 ;
        RECT 40.060 -8.370 40.230 -7.500 ;
        RECT 40.610 -8.370 40.780 -7.680 ;
        RECT 44.750 -7.720 44.920 -7.030 ;
        RECT 45.290 -7.890 45.460 -7.020 ;
        RECT 45.730 -7.060 46.150 -6.780 ;
        RECT 47.370 -6.890 47.540 -6.290 ;
        RECT 49.020 -6.380 49.190 -5.500 ;
        RECT 49.360 -5.560 49.650 -5.500 ;
        RECT 50.880 -5.670 51.300 -5.330 ;
        RECT 51.560 -5.370 51.730 -4.500 ;
        RECT 52.110 -5.370 52.280 -4.680 ;
        RECT 56.250 -4.720 56.420 -4.030 ;
        RECT 56.790 -4.890 56.960 -4.020 ;
        RECT 57.230 -4.060 57.650 -3.780 ;
        RECT 58.870 -3.890 59.040 -3.560 ;
        RECT 60.490 -3.850 60.750 -3.760 ;
        RECT 61.400 -3.850 61.660 -3.760 ;
        RECT 58.170 -4.060 59.590 -3.890 ;
        RECT 60.400 -4.060 60.820 -3.850 ;
        RECT 61.330 -4.060 61.750 -3.850 ;
        RECT 57.230 -4.500 58.810 -4.330 ;
        RECT 60.020 -4.450 60.190 -4.120 ;
        RECT 54.060 -5.270 54.230 -4.940 ;
        RECT 55.470 -5.060 57.050 -4.890 ;
        RECT 52.530 -5.540 52.950 -5.330 ;
        RECT 53.420 -5.540 53.840 -5.330 ;
        RECT 54.650 -5.500 56.110 -5.330 ;
        RECT 52.600 -5.600 52.860 -5.540 ;
        RECT 53.510 -5.600 53.770 -5.540 ;
        RECT 51.020 -6.380 51.190 -5.670 ;
        RECT 48.990 -6.850 49.250 -6.760 ;
        RECT 49.900 -6.850 50.160 -6.760 ;
        RECT 46.670 -7.060 48.090 -6.890 ;
        RECT 48.900 -7.060 49.320 -6.850 ;
        RECT 49.830 -7.060 50.250 -6.850 ;
        RECT 45.730 -7.500 47.310 -7.330 ;
        RECT 48.520 -7.450 48.690 -7.120 ;
        RECT 42.560 -8.270 42.730 -7.940 ;
        RECT 43.970 -8.060 45.550 -7.890 ;
        RECT 41.030 -8.540 41.450 -8.330 ;
        RECT 41.920 -8.540 42.340 -8.330 ;
        RECT 43.150 -8.500 44.610 -8.330 ;
        RECT 41.100 -8.600 41.360 -8.540 ;
        RECT 42.010 -8.600 42.270 -8.540 ;
        RECT 43.610 -8.560 43.900 -8.500 ;
        RECT 45.130 -8.670 45.550 -8.330 ;
        RECT 45.810 -8.370 45.980 -7.500 ;
        RECT 46.360 -8.370 46.530 -7.680 ;
        RECT 50.500 -7.720 50.670 -7.030 ;
        RECT 51.040 -7.890 51.210 -7.020 ;
        RECT 51.480 -7.060 51.900 -6.780 ;
        RECT 53.120 -6.890 53.290 -6.290 ;
        RECT 54.770 -6.380 54.940 -5.500 ;
        RECT 55.110 -5.560 55.400 -5.500 ;
        RECT 56.630 -5.670 57.050 -5.330 ;
        RECT 57.310 -5.370 57.480 -4.500 ;
        RECT 57.860 -5.370 58.030 -4.680 ;
        RECT 62.000 -4.720 62.170 -4.030 ;
        RECT 62.540 -4.890 62.710 -4.020 ;
        RECT 62.980 -4.060 63.400 -3.780 ;
        RECT 64.620 -3.890 64.790 -3.560 ;
        RECT 66.240 -3.850 66.500 -3.760 ;
        RECT 67.150 -3.850 67.410 -3.760 ;
        RECT 63.920 -4.060 65.340 -3.890 ;
        RECT 66.150 -4.060 66.570 -3.850 ;
        RECT 67.080 -4.060 67.500 -3.850 ;
        RECT 62.980 -4.500 64.560 -4.330 ;
        RECT 65.770 -4.450 65.940 -4.120 ;
        RECT 59.810 -5.270 59.980 -4.940 ;
        RECT 61.220 -5.060 62.800 -4.890 ;
        RECT 58.280 -5.540 58.700 -5.330 ;
        RECT 59.170 -5.540 59.590 -5.330 ;
        RECT 60.400 -5.500 61.860 -5.330 ;
        RECT 58.350 -5.600 58.610 -5.540 ;
        RECT 59.260 -5.600 59.520 -5.540 ;
        RECT 56.770 -6.380 56.940 -5.670 ;
        RECT 54.740 -6.850 55.000 -6.760 ;
        RECT 55.650 -6.850 55.910 -6.760 ;
        RECT 52.420 -7.060 53.840 -6.890 ;
        RECT 54.650 -7.060 55.070 -6.850 ;
        RECT 55.580 -7.060 56.000 -6.850 ;
        RECT 51.480 -7.500 53.060 -7.330 ;
        RECT 54.270 -7.450 54.440 -7.120 ;
        RECT 48.310 -8.270 48.480 -7.940 ;
        RECT 49.720 -8.060 51.300 -7.890 ;
        RECT 46.780 -8.540 47.200 -8.330 ;
        RECT 47.670 -8.540 48.090 -8.330 ;
        RECT 48.900 -8.500 50.360 -8.330 ;
        RECT 46.850 -8.600 47.110 -8.540 ;
        RECT 47.760 -8.600 48.020 -8.540 ;
        RECT 49.360 -8.560 49.650 -8.500 ;
        RECT 50.880 -8.670 51.300 -8.330 ;
        RECT 51.560 -8.370 51.730 -7.500 ;
        RECT 52.110 -8.370 52.280 -7.680 ;
        RECT 56.250 -7.720 56.420 -7.030 ;
        RECT 56.790 -7.890 56.960 -7.020 ;
        RECT 57.230 -7.060 57.650 -6.780 ;
        RECT 58.870 -6.890 59.040 -6.290 ;
        RECT 60.520 -6.380 60.690 -5.500 ;
        RECT 60.860 -5.560 61.150 -5.500 ;
        RECT 62.380 -5.670 62.800 -5.330 ;
        RECT 63.060 -5.370 63.230 -4.500 ;
        RECT 63.610 -5.370 63.780 -4.680 ;
        RECT 67.750 -4.720 67.920 -4.030 ;
        RECT 68.290 -4.890 68.460 -4.020 ;
        RECT 68.730 -4.060 69.150 -3.780 ;
        RECT 70.370 -3.890 70.540 -3.560 ;
        RECT 71.990 -3.850 72.250 -3.760 ;
        RECT 72.900 -3.850 73.160 -3.760 ;
        RECT 69.670 -4.060 71.090 -3.890 ;
        RECT 71.900 -4.060 72.320 -3.850 ;
        RECT 72.830 -4.060 73.250 -3.850 ;
        RECT 68.730 -4.500 70.310 -4.330 ;
        RECT 71.520 -4.450 71.690 -4.120 ;
        RECT 65.560 -5.270 65.730 -4.940 ;
        RECT 66.970 -5.060 68.550 -4.890 ;
        RECT 64.030 -5.540 64.450 -5.330 ;
        RECT 64.920 -5.540 65.340 -5.330 ;
        RECT 66.150 -5.500 67.610 -5.330 ;
        RECT 64.100 -5.600 64.360 -5.540 ;
        RECT 65.010 -5.600 65.270 -5.540 ;
        RECT 62.520 -6.380 62.690 -5.670 ;
        RECT 60.490 -6.850 60.750 -6.760 ;
        RECT 61.400 -6.850 61.660 -6.760 ;
        RECT 58.170 -7.060 59.590 -6.890 ;
        RECT 60.400 -7.060 60.820 -6.850 ;
        RECT 61.330 -7.060 61.750 -6.850 ;
        RECT 57.230 -7.500 58.810 -7.330 ;
        RECT 60.020 -7.450 60.190 -7.120 ;
        RECT 54.060 -8.270 54.230 -7.940 ;
        RECT 55.470 -8.060 57.050 -7.890 ;
        RECT 52.530 -8.540 52.950 -8.330 ;
        RECT 53.420 -8.540 53.840 -8.330 ;
        RECT 54.650 -8.500 56.110 -8.330 ;
        RECT 52.600 -8.600 52.860 -8.540 ;
        RECT 53.510 -8.600 53.770 -8.540 ;
        RECT 55.110 -8.560 55.400 -8.500 ;
        RECT 56.630 -8.670 57.050 -8.330 ;
        RECT 57.310 -8.370 57.480 -7.500 ;
        RECT 57.860 -8.370 58.030 -7.680 ;
        RECT 62.000 -7.720 62.170 -7.030 ;
        RECT 62.540 -7.890 62.710 -7.020 ;
        RECT 62.980 -7.060 63.400 -6.780 ;
        RECT 64.620 -6.890 64.790 -6.290 ;
        RECT 66.270 -6.380 66.440 -5.500 ;
        RECT 66.610 -5.560 66.900 -5.500 ;
        RECT 68.130 -5.670 68.550 -5.330 ;
        RECT 68.810 -5.370 68.980 -4.500 ;
        RECT 69.360 -5.370 69.530 -4.680 ;
        RECT 73.500 -4.720 73.670 -4.030 ;
        RECT 74.040 -4.890 74.210 -4.020 ;
        RECT 74.480 -4.060 74.900 -3.780 ;
        RECT 76.120 -3.890 76.290 -3.560 ;
        RECT 77.740 -3.850 78.000 -3.760 ;
        RECT 78.650 -3.850 78.910 -3.760 ;
        RECT 75.420 -4.060 76.840 -3.890 ;
        RECT 77.650 -4.060 78.070 -3.850 ;
        RECT 78.580 -4.060 79.000 -3.850 ;
        RECT 74.480 -4.500 76.060 -4.330 ;
        RECT 77.270 -4.450 77.440 -4.120 ;
        RECT 71.310 -5.270 71.480 -4.940 ;
        RECT 72.720 -5.060 74.300 -4.890 ;
        RECT 69.780 -5.540 70.200 -5.330 ;
        RECT 70.670 -5.540 71.090 -5.330 ;
        RECT 71.900 -5.500 73.360 -5.330 ;
        RECT 69.850 -5.600 70.110 -5.540 ;
        RECT 70.760 -5.600 71.020 -5.540 ;
        RECT 68.270 -6.380 68.440 -5.670 ;
        RECT 66.240 -6.850 66.500 -6.760 ;
        RECT 67.150 -6.850 67.410 -6.760 ;
        RECT 63.920 -7.060 65.340 -6.890 ;
        RECT 66.150 -7.060 66.570 -6.850 ;
        RECT 67.080 -7.060 67.500 -6.850 ;
        RECT 62.980 -7.500 64.560 -7.330 ;
        RECT 65.770 -7.450 65.940 -7.120 ;
        RECT 59.810 -8.270 59.980 -7.940 ;
        RECT 61.220 -8.060 62.800 -7.890 ;
        RECT 58.280 -8.540 58.700 -8.330 ;
        RECT 59.170 -8.540 59.590 -8.330 ;
        RECT 60.400 -8.500 61.860 -8.330 ;
        RECT 58.350 -8.600 58.610 -8.540 ;
        RECT 59.260 -8.600 59.520 -8.540 ;
        RECT 60.860 -8.560 61.150 -8.500 ;
        RECT 62.380 -8.670 62.800 -8.330 ;
        RECT 63.060 -8.370 63.230 -7.500 ;
        RECT 63.610 -8.370 63.780 -7.680 ;
        RECT 67.750 -7.720 67.920 -7.030 ;
        RECT 68.290 -7.890 68.460 -7.020 ;
        RECT 68.730 -7.060 69.150 -6.780 ;
        RECT 70.370 -6.890 70.540 -6.290 ;
        RECT 72.020 -6.380 72.190 -5.500 ;
        RECT 72.360 -5.560 72.650 -5.500 ;
        RECT 73.880 -5.670 74.300 -5.330 ;
        RECT 74.560 -5.370 74.730 -4.500 ;
        RECT 75.110 -5.370 75.280 -4.680 ;
        RECT 79.250 -4.720 79.420 -4.030 ;
        RECT 79.790 -4.890 79.960 -4.020 ;
        RECT 80.230 -4.060 80.650 -3.780 ;
        RECT 81.870 -3.890 82.040 -3.560 ;
        RECT 83.490 -3.850 83.750 -3.760 ;
        RECT 84.400 -3.850 84.660 -3.760 ;
        RECT 81.170 -4.060 82.590 -3.890 ;
        RECT 83.400 -4.060 83.820 -3.850 ;
        RECT 84.330 -4.060 84.750 -3.850 ;
        RECT 80.230 -4.500 81.810 -4.330 ;
        RECT 83.020 -4.450 83.190 -4.120 ;
        RECT 77.060 -5.270 77.230 -4.940 ;
        RECT 78.470 -5.060 80.050 -4.890 ;
        RECT 75.530 -5.540 75.950 -5.330 ;
        RECT 76.420 -5.540 76.840 -5.330 ;
        RECT 77.650 -5.500 79.110 -5.330 ;
        RECT 75.600 -5.600 75.860 -5.540 ;
        RECT 76.510 -5.600 76.770 -5.540 ;
        RECT 74.020 -6.380 74.190 -5.670 ;
        RECT 71.990 -6.850 72.250 -6.760 ;
        RECT 72.900 -6.850 73.160 -6.760 ;
        RECT 69.670 -7.060 71.090 -6.890 ;
        RECT 71.900 -7.060 72.320 -6.850 ;
        RECT 72.830 -7.060 73.250 -6.850 ;
        RECT 68.730 -7.500 70.310 -7.330 ;
        RECT 71.520 -7.450 71.690 -7.120 ;
        RECT 65.560 -8.270 65.730 -7.940 ;
        RECT 66.970 -8.060 68.550 -7.890 ;
        RECT 64.030 -8.540 64.450 -8.330 ;
        RECT 64.920 -8.540 65.340 -8.330 ;
        RECT 66.150 -8.500 67.610 -8.330 ;
        RECT 64.100 -8.600 64.360 -8.540 ;
        RECT 65.010 -8.600 65.270 -8.540 ;
        RECT 66.610 -8.560 66.900 -8.500 ;
        RECT 68.130 -8.670 68.550 -8.330 ;
        RECT 68.810 -8.370 68.980 -7.500 ;
        RECT 69.360 -8.370 69.530 -7.680 ;
        RECT 73.500 -7.720 73.670 -7.030 ;
        RECT 74.040 -7.890 74.210 -7.020 ;
        RECT 74.480 -7.060 74.900 -6.780 ;
        RECT 76.120 -6.890 76.290 -6.290 ;
        RECT 77.770 -6.380 77.940 -5.500 ;
        RECT 78.110 -5.560 78.400 -5.500 ;
        RECT 79.630 -5.670 80.050 -5.330 ;
        RECT 80.310 -5.370 80.480 -4.500 ;
        RECT 80.860 -5.370 81.030 -4.680 ;
        RECT 85.000 -4.720 85.170 -4.030 ;
        RECT 85.540 -4.890 85.710 -4.020 ;
        RECT 85.980 -4.060 86.400 -3.780 ;
        RECT 87.620 -3.890 87.790 -3.560 ;
        RECT 89.240 -3.850 89.500 -3.760 ;
        RECT 90.150 -3.850 90.410 -3.760 ;
        RECT 86.920 -4.060 88.340 -3.890 ;
        RECT 89.150 -4.060 89.570 -3.850 ;
        RECT 90.080 -4.060 90.500 -3.850 ;
        RECT 85.980 -4.500 87.560 -4.330 ;
        RECT 88.770 -4.450 88.940 -4.120 ;
        RECT 82.810 -5.270 82.980 -4.940 ;
        RECT 84.220 -5.060 85.800 -4.890 ;
        RECT 81.280 -5.540 81.700 -5.330 ;
        RECT 82.170 -5.540 82.590 -5.330 ;
        RECT 83.400 -5.500 84.860 -5.330 ;
        RECT 81.350 -5.600 81.610 -5.540 ;
        RECT 82.260 -5.600 82.520 -5.540 ;
        RECT 79.770 -6.380 79.940 -5.670 ;
        RECT 77.740 -6.850 78.000 -6.760 ;
        RECT 78.650 -6.850 78.910 -6.760 ;
        RECT 75.420 -7.060 76.840 -6.890 ;
        RECT 77.650 -7.060 78.070 -6.850 ;
        RECT 78.580 -7.060 79.000 -6.850 ;
        RECT 74.480 -7.500 76.060 -7.330 ;
        RECT 77.270 -7.450 77.440 -7.120 ;
        RECT 71.310 -8.270 71.480 -7.940 ;
        RECT 72.720 -8.060 74.300 -7.890 ;
        RECT 69.780 -8.540 70.200 -8.330 ;
        RECT 70.670 -8.540 71.090 -8.330 ;
        RECT 71.900 -8.500 73.360 -8.330 ;
        RECT 69.850 -8.600 70.110 -8.540 ;
        RECT 70.760 -8.600 71.020 -8.540 ;
        RECT 72.360 -8.560 72.650 -8.500 ;
        RECT 73.880 -8.670 74.300 -8.330 ;
        RECT 74.560 -8.370 74.730 -7.500 ;
        RECT 75.110 -8.370 75.280 -7.680 ;
        RECT 79.250 -7.720 79.420 -7.030 ;
        RECT 79.790 -7.890 79.960 -7.020 ;
        RECT 80.230 -7.060 80.650 -6.780 ;
        RECT 81.870 -6.890 82.040 -6.290 ;
        RECT 83.520 -6.380 83.690 -5.500 ;
        RECT 83.860 -5.560 84.150 -5.500 ;
        RECT 85.380 -5.670 85.800 -5.330 ;
        RECT 86.060 -5.370 86.230 -4.500 ;
        RECT 86.610 -5.370 86.780 -4.680 ;
        RECT 90.750 -4.720 90.920 -4.030 ;
        RECT 91.290 -4.890 91.460 -4.020 ;
        RECT 91.730 -4.060 92.150 -3.780 ;
        RECT 93.370 -3.890 93.540 -3.560 ;
        RECT 92.670 -4.060 94.090 -3.890 ;
        RECT 91.730 -4.500 93.310 -4.330 ;
        RECT 88.560 -5.270 88.730 -4.940 ;
        RECT 89.970 -5.060 91.550 -4.890 ;
        RECT 87.030 -5.540 87.450 -5.330 ;
        RECT 87.920 -5.540 88.340 -5.330 ;
        RECT 89.150 -5.500 90.610 -5.330 ;
        RECT 87.100 -5.600 87.360 -5.540 ;
        RECT 88.010 -5.600 88.270 -5.540 ;
        RECT 85.520 -6.380 85.690 -5.670 ;
        RECT 83.490 -6.850 83.750 -6.760 ;
        RECT 84.400 -6.850 84.660 -6.760 ;
        RECT 81.170 -7.060 82.590 -6.890 ;
        RECT 83.400 -7.060 83.820 -6.850 ;
        RECT 84.330 -7.060 84.750 -6.850 ;
        RECT 80.230 -7.500 81.810 -7.330 ;
        RECT 83.020 -7.450 83.190 -7.120 ;
        RECT 77.060 -8.270 77.230 -7.940 ;
        RECT 78.470 -8.060 80.050 -7.890 ;
        RECT 75.530 -8.540 75.950 -8.330 ;
        RECT 76.420 -8.540 76.840 -8.330 ;
        RECT 77.650 -8.500 79.110 -8.330 ;
        RECT 75.600 -8.600 75.860 -8.540 ;
        RECT 76.510 -8.600 76.770 -8.540 ;
        RECT 78.110 -8.560 78.400 -8.500 ;
        RECT 79.630 -8.670 80.050 -8.330 ;
        RECT 80.310 -8.370 80.480 -7.500 ;
        RECT 80.860 -8.370 81.030 -7.680 ;
        RECT 85.000 -7.720 85.170 -7.030 ;
        RECT 85.540 -7.890 85.710 -7.020 ;
        RECT 85.980 -7.060 86.400 -6.780 ;
        RECT 87.620 -6.890 87.790 -6.290 ;
        RECT 89.270 -6.380 89.440 -5.500 ;
        RECT 89.610 -5.560 89.900 -5.500 ;
        RECT 91.130 -5.670 91.550 -5.330 ;
        RECT 91.810 -5.370 91.980 -4.500 ;
        RECT 92.360 -5.370 92.530 -4.680 ;
        RECT 94.310 -5.270 94.480 -4.940 ;
        RECT 92.780 -5.540 93.200 -5.330 ;
        RECT 93.670 -5.540 94.090 -5.330 ;
        RECT 92.850 -5.600 93.110 -5.540 ;
        RECT 93.760 -5.600 94.020 -5.540 ;
        RECT 91.270 -6.380 91.440 -5.670 ;
        RECT 94.230 -6.290 94.400 -6.020 ;
        RECT 93.370 -6.460 94.400 -6.290 ;
        RECT 89.240 -6.850 89.500 -6.760 ;
        RECT 90.150 -6.850 90.410 -6.760 ;
        RECT 86.920 -7.060 88.340 -6.890 ;
        RECT 89.150 -7.060 89.570 -6.850 ;
        RECT 90.080 -7.060 90.500 -6.850 ;
        RECT 85.980 -7.500 87.560 -7.330 ;
        RECT 88.770 -7.450 88.940 -7.120 ;
        RECT 82.810 -8.270 82.980 -7.940 ;
        RECT 84.220 -8.060 85.800 -7.890 ;
        RECT 81.280 -8.540 81.700 -8.330 ;
        RECT 82.170 -8.540 82.590 -8.330 ;
        RECT 83.400 -8.500 84.860 -8.330 ;
        RECT 81.350 -8.600 81.610 -8.540 ;
        RECT 82.260 -8.600 82.520 -8.540 ;
        RECT 83.860 -8.560 84.150 -8.500 ;
        RECT 85.380 -8.670 85.800 -8.330 ;
        RECT 86.060 -8.370 86.230 -7.500 ;
        RECT 86.610 -8.370 86.780 -7.680 ;
        RECT 90.750 -7.720 90.920 -7.030 ;
        RECT 91.290 -7.890 91.460 -7.020 ;
        RECT 91.730 -7.060 92.150 -6.780 ;
        RECT 93.370 -6.890 93.540 -6.460 ;
        RECT 92.670 -7.060 94.090 -6.890 ;
        RECT 91.730 -7.500 93.310 -7.330 ;
        RECT 88.560 -8.270 88.730 -7.940 ;
        RECT 89.970 -8.060 91.550 -7.890 ;
        RECT 87.030 -8.540 87.450 -8.330 ;
        RECT 87.920 -8.540 88.340 -8.330 ;
        RECT 89.150 -8.500 90.610 -8.330 ;
        RECT 87.100 -8.600 87.360 -8.540 ;
        RECT 88.010 -8.600 88.270 -8.540 ;
        RECT 89.610 -8.560 89.900 -8.500 ;
        RECT 91.130 -8.670 91.550 -8.330 ;
        RECT 91.810 -8.370 91.980 -7.500 ;
        RECT 92.360 -8.370 92.530 -7.680 ;
        RECT 94.310 -8.270 94.480 -7.940 ;
        RECT 92.780 -8.540 93.200 -8.330 ;
        RECT 93.670 -8.540 94.090 -8.330 ;
        RECT 92.850 -8.600 93.110 -8.540 ;
        RECT 93.760 -8.600 94.020 -8.540 ;
        RECT 2.990 -9.260 3.250 -9.170 ;
        RECT 3.900 -9.260 4.160 -9.170 ;
        RECT 2.900 -9.470 3.320 -9.260 ;
        RECT 3.830 -9.470 4.250 -9.260 ;
        RECT 2.520 -9.860 2.690 -9.530 ;
        RECT 4.500 -10.130 4.670 -9.440 ;
        RECT 5.040 -10.300 5.210 -9.430 ;
        RECT 5.480 -9.470 5.900 -9.190 ;
        RECT 7.120 -9.300 7.290 -8.970 ;
        RECT 8.740 -9.260 9.000 -9.170 ;
        RECT 9.650 -9.260 9.910 -9.170 ;
        RECT 6.420 -9.470 7.840 -9.300 ;
        RECT 8.650 -9.470 9.070 -9.260 ;
        RECT 9.580 -9.470 10.000 -9.260 ;
        RECT 5.480 -9.910 7.060 -9.740 ;
        RECT 8.270 -9.860 8.440 -9.530 ;
        RECT 3.720 -10.470 5.300 -10.300 ;
        RECT 2.900 -10.910 4.360 -10.740 ;
        RECT 3.360 -10.970 3.650 -10.910 ;
        RECT 4.880 -11.080 5.300 -10.740 ;
        RECT 5.560 -10.780 5.730 -9.910 ;
        RECT 6.110 -10.780 6.280 -10.090 ;
        RECT 10.250 -10.130 10.420 -9.440 ;
        RECT 10.790 -10.300 10.960 -9.430 ;
        RECT 11.230 -9.470 11.650 -9.190 ;
        RECT 12.870 -9.300 13.040 -8.970 ;
        RECT 14.490 -9.260 14.750 -9.170 ;
        RECT 15.400 -9.260 15.660 -9.170 ;
        RECT 12.170 -9.470 13.590 -9.300 ;
        RECT 14.400 -9.470 14.820 -9.260 ;
        RECT 15.330 -9.470 15.750 -9.260 ;
        RECT 11.230 -9.910 12.810 -9.740 ;
        RECT 14.020 -9.860 14.190 -9.530 ;
        RECT 8.060 -10.680 8.230 -10.350 ;
        RECT 9.470 -10.470 11.050 -10.300 ;
        RECT 6.530 -10.950 6.950 -10.740 ;
        RECT 7.420 -10.950 7.840 -10.740 ;
        RECT 8.650 -10.910 10.110 -10.740 ;
        RECT 6.600 -11.010 6.860 -10.950 ;
        RECT 7.510 -11.010 7.770 -10.950 ;
        RECT 9.110 -10.970 9.400 -10.910 ;
        RECT 10.630 -11.080 11.050 -10.740 ;
        RECT 11.310 -10.780 11.480 -9.910 ;
        RECT 11.860 -10.780 12.030 -10.090 ;
        RECT 16.000 -10.130 16.170 -9.440 ;
        RECT 16.540 -10.300 16.710 -9.430 ;
        RECT 16.980 -9.470 17.400 -9.190 ;
        RECT 18.620 -9.300 18.790 -8.970 ;
        RECT 20.240 -9.260 20.500 -9.170 ;
        RECT 21.150 -9.260 21.410 -9.170 ;
        RECT 17.920 -9.470 19.340 -9.300 ;
        RECT 20.150 -9.470 20.570 -9.260 ;
        RECT 21.080 -9.470 21.500 -9.260 ;
        RECT 16.980 -9.910 18.560 -9.740 ;
        RECT 19.770 -9.860 19.940 -9.530 ;
        RECT 13.810 -10.680 13.980 -10.350 ;
        RECT 15.220 -10.470 16.800 -10.300 ;
        RECT 12.280 -10.950 12.700 -10.740 ;
        RECT 13.170 -10.950 13.590 -10.740 ;
        RECT 14.400 -10.910 15.860 -10.740 ;
        RECT 12.350 -11.010 12.610 -10.950 ;
        RECT 13.260 -11.010 13.520 -10.950 ;
        RECT 14.860 -10.970 15.150 -10.910 ;
        RECT 16.380 -11.080 16.800 -10.740 ;
        RECT 17.060 -10.780 17.230 -9.910 ;
        RECT 17.610 -10.780 17.780 -10.090 ;
        RECT 21.750 -10.130 21.920 -9.440 ;
        RECT 22.290 -10.300 22.460 -9.430 ;
        RECT 22.730 -9.470 23.150 -9.190 ;
        RECT 24.370 -9.300 24.540 -8.970 ;
        RECT 25.990 -9.260 26.250 -9.170 ;
        RECT 26.900 -9.260 27.160 -9.170 ;
        RECT 23.670 -9.470 25.090 -9.300 ;
        RECT 25.900 -9.470 26.320 -9.260 ;
        RECT 26.830 -9.470 27.250 -9.260 ;
        RECT 22.730 -9.910 24.310 -9.740 ;
        RECT 25.520 -9.860 25.690 -9.530 ;
        RECT 19.560 -10.680 19.730 -10.350 ;
        RECT 20.970 -10.470 22.550 -10.300 ;
        RECT 18.030 -10.950 18.450 -10.740 ;
        RECT 18.920 -10.950 19.340 -10.740 ;
        RECT 20.150 -10.910 21.610 -10.740 ;
        RECT 18.100 -11.010 18.360 -10.950 ;
        RECT 19.010 -11.010 19.270 -10.950 ;
        RECT 20.610 -10.970 20.900 -10.910 ;
        RECT 22.130 -11.080 22.550 -10.740 ;
        RECT 22.810 -10.780 22.980 -9.910 ;
        RECT 23.360 -10.780 23.530 -10.090 ;
        RECT 27.500 -10.130 27.670 -9.440 ;
        RECT 28.040 -10.300 28.210 -9.430 ;
        RECT 28.480 -9.470 28.900 -9.190 ;
        RECT 30.120 -9.300 30.290 -8.970 ;
        RECT 31.740 -9.260 32.000 -9.170 ;
        RECT 32.650 -9.260 32.910 -9.170 ;
        RECT 29.420 -9.470 30.840 -9.300 ;
        RECT 31.650 -9.470 32.070 -9.260 ;
        RECT 32.580 -9.470 33.000 -9.260 ;
        RECT 28.480 -9.910 30.060 -9.740 ;
        RECT 31.270 -9.860 31.440 -9.530 ;
        RECT 25.310 -10.680 25.480 -10.350 ;
        RECT 26.720 -10.470 28.300 -10.300 ;
        RECT 23.780 -10.950 24.200 -10.740 ;
        RECT 24.670 -10.950 25.090 -10.740 ;
        RECT 25.900 -10.910 27.360 -10.740 ;
        RECT 23.850 -11.010 24.110 -10.950 ;
        RECT 24.760 -11.010 25.020 -10.950 ;
        RECT 26.360 -10.970 26.650 -10.910 ;
        RECT 27.880 -11.080 28.300 -10.740 ;
        RECT 28.560 -10.780 28.730 -9.910 ;
        RECT 29.110 -10.780 29.280 -10.090 ;
        RECT 33.250 -10.130 33.420 -9.440 ;
        RECT 33.790 -10.300 33.960 -9.430 ;
        RECT 34.230 -9.470 34.650 -9.190 ;
        RECT 35.870 -9.300 36.040 -8.970 ;
        RECT 37.490 -9.260 37.750 -9.170 ;
        RECT 38.400 -9.260 38.660 -9.170 ;
        RECT 35.170 -9.470 36.590 -9.300 ;
        RECT 37.400 -9.470 37.820 -9.260 ;
        RECT 38.330 -9.470 38.750 -9.260 ;
        RECT 34.230 -9.910 35.810 -9.740 ;
        RECT 37.020 -9.860 37.190 -9.530 ;
        RECT 31.060 -10.680 31.230 -10.350 ;
        RECT 32.470 -10.470 34.050 -10.300 ;
        RECT 29.530 -10.950 29.950 -10.740 ;
        RECT 30.420 -10.950 30.840 -10.740 ;
        RECT 31.650 -10.910 33.110 -10.740 ;
        RECT 29.600 -11.010 29.860 -10.950 ;
        RECT 30.510 -11.010 30.770 -10.950 ;
        RECT 32.110 -10.970 32.400 -10.910 ;
        RECT 33.630 -11.080 34.050 -10.740 ;
        RECT 34.310 -10.780 34.480 -9.910 ;
        RECT 34.860 -10.780 35.030 -10.090 ;
        RECT 39.000 -10.130 39.170 -9.440 ;
        RECT 39.540 -10.300 39.710 -9.430 ;
        RECT 39.980 -9.470 40.400 -9.190 ;
        RECT 41.620 -9.300 41.790 -8.970 ;
        RECT 43.240 -9.260 43.500 -9.170 ;
        RECT 44.150 -9.260 44.410 -9.170 ;
        RECT 40.920 -9.470 42.340 -9.300 ;
        RECT 43.150 -9.470 43.570 -9.260 ;
        RECT 44.080 -9.470 44.500 -9.260 ;
        RECT 39.980 -9.910 41.560 -9.740 ;
        RECT 42.770 -9.860 42.940 -9.530 ;
        RECT 36.810 -10.680 36.980 -10.350 ;
        RECT 38.220 -10.470 39.800 -10.300 ;
        RECT 35.280 -10.950 35.700 -10.740 ;
        RECT 36.170 -10.950 36.590 -10.740 ;
        RECT 37.400 -10.910 38.860 -10.740 ;
        RECT 35.350 -11.010 35.610 -10.950 ;
        RECT 36.260 -11.010 36.520 -10.950 ;
        RECT 37.860 -10.970 38.150 -10.910 ;
        RECT 39.380 -11.080 39.800 -10.740 ;
        RECT 40.060 -10.780 40.230 -9.910 ;
        RECT 40.610 -10.780 40.780 -10.090 ;
        RECT 44.750 -10.130 44.920 -9.440 ;
        RECT 45.290 -10.300 45.460 -9.430 ;
        RECT 45.730 -9.470 46.150 -9.190 ;
        RECT 47.370 -9.300 47.540 -8.970 ;
        RECT 48.990 -9.260 49.250 -9.170 ;
        RECT 49.900 -9.260 50.160 -9.170 ;
        RECT 46.670 -9.470 48.090 -9.300 ;
        RECT 48.900 -9.470 49.320 -9.260 ;
        RECT 49.830 -9.470 50.250 -9.260 ;
        RECT 45.730 -9.910 47.310 -9.740 ;
        RECT 48.520 -9.860 48.690 -9.530 ;
        RECT 42.560 -10.680 42.730 -10.350 ;
        RECT 43.970 -10.470 45.550 -10.300 ;
        RECT 41.030 -10.950 41.450 -10.740 ;
        RECT 41.920 -10.950 42.340 -10.740 ;
        RECT 43.150 -10.910 44.610 -10.740 ;
        RECT 41.100 -11.010 41.360 -10.950 ;
        RECT 42.010 -11.010 42.270 -10.950 ;
        RECT 43.610 -10.970 43.900 -10.910 ;
        RECT 45.130 -11.080 45.550 -10.740 ;
        RECT 45.810 -10.780 45.980 -9.910 ;
        RECT 46.360 -10.780 46.530 -10.090 ;
        RECT 50.500 -10.130 50.670 -9.440 ;
        RECT 51.040 -10.300 51.210 -9.430 ;
        RECT 51.480 -9.470 51.900 -9.190 ;
        RECT 53.120 -9.300 53.290 -8.970 ;
        RECT 54.740 -9.260 55.000 -9.170 ;
        RECT 55.650 -9.260 55.910 -9.170 ;
        RECT 52.420 -9.470 53.840 -9.300 ;
        RECT 54.650 -9.470 55.070 -9.260 ;
        RECT 55.580 -9.470 56.000 -9.260 ;
        RECT 51.480 -9.910 53.060 -9.740 ;
        RECT 54.270 -9.860 54.440 -9.530 ;
        RECT 48.310 -10.680 48.480 -10.350 ;
        RECT 49.720 -10.470 51.300 -10.300 ;
        RECT 46.780 -10.950 47.200 -10.740 ;
        RECT 47.670 -10.950 48.090 -10.740 ;
        RECT 48.900 -10.910 50.360 -10.740 ;
        RECT 46.850 -11.010 47.110 -10.950 ;
        RECT 47.760 -11.010 48.020 -10.950 ;
        RECT 49.360 -10.970 49.650 -10.910 ;
        RECT 50.880 -11.080 51.300 -10.740 ;
        RECT 51.560 -10.780 51.730 -9.910 ;
        RECT 52.110 -10.780 52.280 -10.090 ;
        RECT 56.250 -10.130 56.420 -9.440 ;
        RECT 56.790 -10.300 56.960 -9.430 ;
        RECT 57.230 -9.470 57.650 -9.190 ;
        RECT 58.870 -9.300 59.040 -8.970 ;
        RECT 60.490 -9.260 60.750 -9.170 ;
        RECT 61.400 -9.260 61.660 -9.170 ;
        RECT 58.170 -9.470 59.590 -9.300 ;
        RECT 60.400 -9.470 60.820 -9.260 ;
        RECT 61.330 -9.470 61.750 -9.260 ;
        RECT 57.230 -9.910 58.810 -9.740 ;
        RECT 60.020 -9.860 60.190 -9.530 ;
        RECT 54.060 -10.680 54.230 -10.350 ;
        RECT 55.470 -10.470 57.050 -10.300 ;
        RECT 52.530 -10.950 52.950 -10.740 ;
        RECT 53.420 -10.950 53.840 -10.740 ;
        RECT 54.650 -10.910 56.110 -10.740 ;
        RECT 52.600 -11.010 52.860 -10.950 ;
        RECT 53.510 -11.010 53.770 -10.950 ;
        RECT 55.110 -10.970 55.400 -10.910 ;
        RECT 56.630 -11.080 57.050 -10.740 ;
        RECT 57.310 -10.780 57.480 -9.910 ;
        RECT 57.860 -10.780 58.030 -10.090 ;
        RECT 62.000 -10.130 62.170 -9.440 ;
        RECT 62.540 -10.300 62.710 -9.430 ;
        RECT 62.980 -9.470 63.400 -9.190 ;
        RECT 64.620 -9.300 64.790 -8.970 ;
        RECT 66.240 -9.260 66.500 -9.170 ;
        RECT 67.150 -9.260 67.410 -9.170 ;
        RECT 63.920 -9.470 65.340 -9.300 ;
        RECT 66.150 -9.470 66.570 -9.260 ;
        RECT 67.080 -9.470 67.500 -9.260 ;
        RECT 62.980 -9.910 64.560 -9.740 ;
        RECT 65.770 -9.860 65.940 -9.530 ;
        RECT 59.810 -10.680 59.980 -10.350 ;
        RECT 61.220 -10.470 62.800 -10.300 ;
        RECT 58.280 -10.950 58.700 -10.740 ;
        RECT 59.170 -10.950 59.590 -10.740 ;
        RECT 60.400 -10.910 61.860 -10.740 ;
        RECT 58.350 -11.010 58.610 -10.950 ;
        RECT 59.260 -11.010 59.520 -10.950 ;
        RECT 60.860 -10.970 61.150 -10.910 ;
        RECT 62.380 -11.080 62.800 -10.740 ;
        RECT 63.060 -10.780 63.230 -9.910 ;
        RECT 63.610 -10.780 63.780 -10.090 ;
        RECT 67.750 -10.130 67.920 -9.440 ;
        RECT 68.290 -10.300 68.460 -9.430 ;
        RECT 68.730 -9.470 69.150 -9.190 ;
        RECT 70.370 -9.300 70.540 -8.970 ;
        RECT 71.990 -9.260 72.250 -9.170 ;
        RECT 72.900 -9.260 73.160 -9.170 ;
        RECT 69.670 -9.470 71.090 -9.300 ;
        RECT 71.900 -9.470 72.320 -9.260 ;
        RECT 72.830 -9.470 73.250 -9.260 ;
        RECT 68.730 -9.910 70.310 -9.740 ;
        RECT 71.520 -9.860 71.690 -9.530 ;
        RECT 65.560 -10.680 65.730 -10.350 ;
        RECT 66.970 -10.470 68.550 -10.300 ;
        RECT 64.030 -10.950 64.450 -10.740 ;
        RECT 64.920 -10.950 65.340 -10.740 ;
        RECT 66.150 -10.910 67.610 -10.740 ;
        RECT 64.100 -11.010 64.360 -10.950 ;
        RECT 65.010 -11.010 65.270 -10.950 ;
        RECT 66.610 -10.970 66.900 -10.910 ;
        RECT 68.130 -11.080 68.550 -10.740 ;
        RECT 68.810 -10.780 68.980 -9.910 ;
        RECT 69.360 -10.780 69.530 -10.090 ;
        RECT 73.500 -10.130 73.670 -9.440 ;
        RECT 74.040 -10.300 74.210 -9.430 ;
        RECT 74.480 -9.470 74.900 -9.190 ;
        RECT 76.120 -9.300 76.290 -8.970 ;
        RECT 77.740 -9.260 78.000 -9.170 ;
        RECT 78.650 -9.260 78.910 -9.170 ;
        RECT 75.420 -9.470 76.840 -9.300 ;
        RECT 77.650 -9.470 78.070 -9.260 ;
        RECT 78.580 -9.470 79.000 -9.260 ;
        RECT 74.480 -9.910 76.060 -9.740 ;
        RECT 77.270 -9.860 77.440 -9.530 ;
        RECT 71.310 -10.680 71.480 -10.350 ;
        RECT 72.720 -10.470 74.300 -10.300 ;
        RECT 69.780 -10.950 70.200 -10.740 ;
        RECT 70.670 -10.950 71.090 -10.740 ;
        RECT 71.900 -10.910 73.360 -10.740 ;
        RECT 69.850 -11.010 70.110 -10.950 ;
        RECT 70.760 -11.010 71.020 -10.950 ;
        RECT 72.360 -10.970 72.650 -10.910 ;
        RECT 73.880 -11.080 74.300 -10.740 ;
        RECT 74.560 -10.780 74.730 -9.910 ;
        RECT 75.110 -10.780 75.280 -10.090 ;
        RECT 79.250 -10.130 79.420 -9.440 ;
        RECT 79.790 -10.300 79.960 -9.430 ;
        RECT 80.230 -9.470 80.650 -9.190 ;
        RECT 81.870 -9.300 82.040 -8.970 ;
        RECT 83.490 -9.260 83.750 -9.170 ;
        RECT 84.400 -9.260 84.660 -9.170 ;
        RECT 81.170 -9.470 82.590 -9.300 ;
        RECT 83.400 -9.470 83.820 -9.260 ;
        RECT 84.330 -9.470 84.750 -9.260 ;
        RECT 80.230 -9.910 81.810 -9.740 ;
        RECT 83.020 -9.860 83.190 -9.530 ;
        RECT 77.060 -10.680 77.230 -10.350 ;
        RECT 78.470 -10.470 80.050 -10.300 ;
        RECT 75.530 -10.950 75.950 -10.740 ;
        RECT 76.420 -10.950 76.840 -10.740 ;
        RECT 77.650 -10.910 79.110 -10.740 ;
        RECT 75.600 -11.010 75.860 -10.950 ;
        RECT 76.510 -11.010 76.770 -10.950 ;
        RECT 78.110 -10.970 78.400 -10.910 ;
        RECT 79.630 -11.080 80.050 -10.740 ;
        RECT 80.310 -10.780 80.480 -9.910 ;
        RECT 80.860 -10.780 81.030 -10.090 ;
        RECT 85.000 -10.130 85.170 -9.440 ;
        RECT 85.540 -10.300 85.710 -9.430 ;
        RECT 85.980 -9.470 86.400 -9.190 ;
        RECT 87.620 -9.300 87.790 -8.970 ;
        RECT 89.240 -9.260 89.500 -9.170 ;
        RECT 90.150 -9.260 90.410 -9.170 ;
        RECT 86.920 -9.470 88.340 -9.300 ;
        RECT 89.150 -9.470 89.570 -9.260 ;
        RECT 90.080 -9.470 90.500 -9.260 ;
        RECT 85.980 -9.910 87.560 -9.740 ;
        RECT 88.770 -9.860 88.940 -9.530 ;
        RECT 82.810 -10.680 82.980 -10.350 ;
        RECT 84.220 -10.470 85.800 -10.300 ;
        RECT 81.280 -10.950 81.700 -10.740 ;
        RECT 82.170 -10.950 82.590 -10.740 ;
        RECT 83.400 -10.910 84.860 -10.740 ;
        RECT 81.350 -11.010 81.610 -10.950 ;
        RECT 82.260 -11.010 82.520 -10.950 ;
        RECT 83.860 -10.970 84.150 -10.910 ;
        RECT 85.380 -11.080 85.800 -10.740 ;
        RECT 86.060 -10.780 86.230 -9.910 ;
        RECT 86.610 -10.780 86.780 -10.090 ;
        RECT 90.750 -10.130 90.920 -9.440 ;
        RECT 91.290 -10.300 91.460 -9.430 ;
        RECT 91.730 -9.470 92.150 -9.190 ;
        RECT 93.370 -9.300 93.540 -8.970 ;
        RECT 92.670 -9.470 94.090 -9.300 ;
        RECT 91.730 -9.910 93.310 -9.740 ;
        RECT 88.560 -10.680 88.730 -10.350 ;
        RECT 89.970 -10.470 91.550 -10.300 ;
        RECT 87.030 -10.950 87.450 -10.740 ;
        RECT 87.920 -10.950 88.340 -10.740 ;
        RECT 89.150 -10.910 90.610 -10.740 ;
        RECT 87.100 -11.010 87.360 -10.950 ;
        RECT 88.010 -11.010 88.270 -10.950 ;
        RECT 89.610 -10.970 89.900 -10.910 ;
        RECT 91.130 -11.080 91.550 -10.740 ;
        RECT 91.810 -10.780 91.980 -9.910 ;
        RECT 92.360 -10.780 92.530 -10.090 ;
        RECT 94.310 -10.680 94.480 -10.350 ;
        RECT 92.780 -10.950 93.200 -10.740 ;
        RECT 93.670 -10.950 94.090 -10.740 ;
        RECT 92.850 -11.010 93.110 -10.950 ;
        RECT 93.760 -11.010 94.020 -10.950 ;
        RECT 3.140 -13.890 3.310 -11.710 ;
        RECT 3.580 -12.660 3.750 -11.710 ;
        RECT 3.580 -12.830 3.790 -12.660 ;
        RECT 3.580 -13.710 3.750 -12.830 ;
        RECT 4.600 -13.890 4.770 -11.710 ;
        RECT 5.040 -12.660 5.210 -11.710 ;
        RECT 5.570 -12.660 5.740 -11.710 ;
        RECT 5.040 -12.830 5.740 -12.660 ;
        RECT 5.040 -13.710 5.210 -12.830 ;
        RECT 5.570 -13.710 5.740 -12.830 ;
        RECT 3.140 -14.060 4.770 -13.890 ;
        RECT 6.010 -13.890 6.180 -11.710 ;
        RECT 7.000 -12.660 7.170 -11.710 ;
        RECT 6.960 -12.830 7.170 -12.660 ;
        RECT 7.000 -13.710 7.170 -12.830 ;
        RECT 7.440 -13.890 7.610 -11.710 ;
        RECT 6.010 -13.950 7.610 -13.890 ;
        RECT 4.600 -14.290 4.770 -14.060 ;
        RECT 4.950 -14.060 7.610 -13.950 ;
        RECT 8.890 -13.890 9.060 -11.710 ;
        RECT 9.330 -12.660 9.500 -11.710 ;
        RECT 9.330 -12.830 9.540 -12.660 ;
        RECT 9.330 -13.710 9.500 -12.830 ;
        RECT 10.350 -13.890 10.520 -11.710 ;
        RECT 10.790 -12.660 10.960 -11.710 ;
        RECT 11.320 -12.660 11.490 -11.710 ;
        RECT 10.790 -12.830 11.490 -12.660 ;
        RECT 10.790 -13.710 10.960 -12.830 ;
        RECT 11.320 -13.710 11.490 -12.830 ;
        RECT 8.890 -14.060 10.520 -13.890 ;
        RECT 11.760 -13.890 11.930 -11.710 ;
        RECT 12.750 -12.660 12.920 -11.710 ;
        RECT 12.710 -12.830 12.920 -12.660 ;
        RECT 12.750 -13.710 12.920 -12.830 ;
        RECT 13.190 -13.890 13.360 -11.710 ;
        RECT 11.760 -13.950 13.360 -13.890 ;
        RECT 4.950 -14.120 6.180 -14.060 ;
        RECT 3.330 -14.490 3.660 -14.320 ;
        RECT 3.870 -14.490 4.200 -14.320 ;
        RECT 4.600 -14.460 5.840 -14.290 ;
        RECT 3.640 -18.180 3.810 -14.700 ;
        RECT 4.080 -17.700 4.250 -14.700 ;
        RECT 4.600 -17.700 4.770 -14.460 ;
        RECT 5.040 -17.700 5.210 -14.700 ;
        RECT 5.570 -17.700 5.740 -14.700 ;
        RECT 6.010 -17.700 6.180 -14.120 ;
        RECT 10.350 -14.290 10.520 -14.060 ;
        RECT 10.700 -14.060 13.360 -13.950 ;
        RECT 14.640 -13.890 14.810 -11.710 ;
        RECT 15.080 -12.660 15.250 -11.710 ;
        RECT 15.080 -12.830 15.290 -12.660 ;
        RECT 15.080 -13.710 15.250 -12.830 ;
        RECT 16.100 -13.890 16.270 -11.710 ;
        RECT 16.540 -12.660 16.710 -11.710 ;
        RECT 17.070 -12.660 17.240 -11.710 ;
        RECT 16.540 -12.830 17.240 -12.660 ;
        RECT 16.540 -13.710 16.710 -12.830 ;
        RECT 17.070 -13.710 17.240 -12.830 ;
        RECT 14.640 -14.060 16.270 -13.890 ;
        RECT 17.510 -13.890 17.680 -11.710 ;
        RECT 18.500 -12.660 18.670 -11.710 ;
        RECT 18.460 -12.830 18.670 -12.660 ;
        RECT 18.500 -13.710 18.670 -12.830 ;
        RECT 18.940 -13.890 19.110 -11.710 ;
        RECT 17.510 -13.950 19.110 -13.890 ;
        RECT 10.700 -14.120 11.930 -14.060 ;
        RECT 6.580 -14.490 6.910 -14.320 ;
        RECT 7.120 -14.490 7.450 -14.320 ;
        RECT 9.080 -14.490 9.410 -14.320 ;
        RECT 9.620 -14.490 9.950 -14.320 ;
        RECT 10.350 -14.460 11.590 -14.290 ;
        RECT 6.530 -17.700 6.700 -14.700 ;
        RECT 6.970 -18.180 7.140 -14.700 ;
        RECT 3.640 -18.350 7.140 -18.180 ;
        RECT 9.390 -18.180 9.560 -14.700 ;
        RECT 9.830 -17.700 10.000 -14.700 ;
        RECT 10.350 -17.700 10.520 -14.460 ;
        RECT 10.790 -17.700 10.960 -14.700 ;
        RECT 11.320 -17.700 11.490 -14.700 ;
        RECT 11.760 -17.700 11.930 -14.120 ;
        RECT 16.100 -14.290 16.270 -14.060 ;
        RECT 16.450 -14.060 19.110 -13.950 ;
        RECT 20.390 -13.890 20.560 -11.710 ;
        RECT 20.830 -12.660 21.000 -11.710 ;
        RECT 20.830 -12.830 21.040 -12.660 ;
        RECT 20.830 -13.710 21.000 -12.830 ;
        RECT 21.850 -13.890 22.020 -11.710 ;
        RECT 22.290 -12.660 22.460 -11.710 ;
        RECT 22.820 -12.660 22.990 -11.710 ;
        RECT 22.290 -12.830 22.990 -12.660 ;
        RECT 22.290 -13.710 22.460 -12.830 ;
        RECT 22.820 -13.710 22.990 -12.830 ;
        RECT 20.390 -14.060 22.020 -13.890 ;
        RECT 23.260 -13.890 23.430 -11.710 ;
        RECT 24.250 -12.660 24.420 -11.710 ;
        RECT 24.210 -12.830 24.420 -12.660 ;
        RECT 24.250 -13.710 24.420 -12.830 ;
        RECT 24.690 -13.890 24.860 -11.710 ;
        RECT 23.260 -13.950 24.860 -13.890 ;
        RECT 16.450 -14.120 17.680 -14.060 ;
        RECT 12.330 -14.490 12.660 -14.320 ;
        RECT 12.870 -14.490 13.200 -14.320 ;
        RECT 14.830 -14.490 15.160 -14.320 ;
        RECT 15.370 -14.490 15.700 -14.320 ;
        RECT 16.100 -14.460 17.340 -14.290 ;
        RECT 12.280 -17.700 12.450 -14.700 ;
        RECT 12.720 -18.180 12.890 -14.700 ;
        RECT 9.390 -18.350 12.890 -18.180 ;
        RECT 15.140 -18.180 15.310 -14.700 ;
        RECT 15.580 -17.700 15.750 -14.700 ;
        RECT 16.100 -17.700 16.270 -14.460 ;
        RECT 16.540 -17.700 16.710 -14.700 ;
        RECT 17.070 -17.700 17.240 -14.700 ;
        RECT 17.510 -17.700 17.680 -14.120 ;
        RECT 21.850 -14.290 22.020 -14.060 ;
        RECT 22.200 -14.060 24.860 -13.950 ;
        RECT 26.140 -13.890 26.310 -11.710 ;
        RECT 26.580 -12.660 26.750 -11.710 ;
        RECT 26.580 -12.830 26.790 -12.660 ;
        RECT 26.580 -13.710 26.750 -12.830 ;
        RECT 27.600 -13.890 27.770 -11.710 ;
        RECT 28.040 -12.660 28.210 -11.710 ;
        RECT 28.570 -12.660 28.740 -11.710 ;
        RECT 28.040 -12.830 28.740 -12.660 ;
        RECT 28.040 -13.710 28.210 -12.830 ;
        RECT 28.570 -13.710 28.740 -12.830 ;
        RECT 26.140 -14.060 27.770 -13.890 ;
        RECT 29.010 -13.890 29.180 -11.710 ;
        RECT 30.000 -12.660 30.170 -11.710 ;
        RECT 29.960 -12.830 30.170 -12.660 ;
        RECT 30.000 -13.710 30.170 -12.830 ;
        RECT 30.440 -13.890 30.610 -11.710 ;
        RECT 29.010 -13.950 30.610 -13.890 ;
        RECT 22.200 -14.120 23.430 -14.060 ;
        RECT 18.080 -14.490 18.410 -14.320 ;
        RECT 18.620 -14.490 18.950 -14.320 ;
        RECT 20.580 -14.490 20.910 -14.320 ;
        RECT 21.120 -14.490 21.450 -14.320 ;
        RECT 21.850 -14.460 23.090 -14.290 ;
        RECT 18.030 -17.700 18.200 -14.700 ;
        RECT 18.470 -18.180 18.640 -14.700 ;
        RECT 15.140 -18.350 18.640 -18.180 ;
        RECT 20.890 -18.180 21.060 -14.700 ;
        RECT 21.330 -17.700 21.500 -14.700 ;
        RECT 21.850 -17.700 22.020 -14.460 ;
        RECT 22.290 -17.700 22.460 -14.700 ;
        RECT 22.820 -17.700 22.990 -14.700 ;
        RECT 23.260 -17.700 23.430 -14.120 ;
        RECT 27.600 -14.290 27.770 -14.060 ;
        RECT 27.950 -14.060 30.610 -13.950 ;
        RECT 31.890 -13.890 32.060 -11.710 ;
        RECT 32.330 -12.660 32.500 -11.710 ;
        RECT 32.330 -12.830 32.540 -12.660 ;
        RECT 32.330 -13.710 32.500 -12.830 ;
        RECT 33.350 -13.890 33.520 -11.710 ;
        RECT 33.790 -12.660 33.960 -11.710 ;
        RECT 34.320 -12.660 34.490 -11.710 ;
        RECT 33.790 -12.830 34.490 -12.660 ;
        RECT 33.790 -13.710 33.960 -12.830 ;
        RECT 34.320 -13.710 34.490 -12.830 ;
        RECT 31.890 -14.060 33.520 -13.890 ;
        RECT 34.760 -13.890 34.930 -11.710 ;
        RECT 35.750 -12.660 35.920 -11.710 ;
        RECT 35.710 -12.830 35.920 -12.660 ;
        RECT 35.750 -13.710 35.920 -12.830 ;
        RECT 36.190 -13.890 36.360 -11.710 ;
        RECT 34.760 -13.950 36.360 -13.890 ;
        RECT 27.950 -14.120 29.180 -14.060 ;
        RECT 23.830 -14.490 24.160 -14.320 ;
        RECT 24.370 -14.490 24.700 -14.320 ;
        RECT 26.330 -14.490 26.660 -14.320 ;
        RECT 26.870 -14.490 27.200 -14.320 ;
        RECT 27.600 -14.460 28.840 -14.290 ;
        RECT 23.780 -17.700 23.950 -14.700 ;
        RECT 24.220 -18.180 24.390 -14.700 ;
        RECT 20.890 -18.350 24.390 -18.180 ;
        RECT 26.640 -18.180 26.810 -14.700 ;
        RECT 27.080 -17.700 27.250 -14.700 ;
        RECT 27.600 -17.700 27.770 -14.460 ;
        RECT 28.040 -17.700 28.210 -14.700 ;
        RECT 28.570 -17.700 28.740 -14.700 ;
        RECT 29.010 -17.700 29.180 -14.120 ;
        RECT 33.350 -14.290 33.520 -14.060 ;
        RECT 33.700 -14.060 36.360 -13.950 ;
        RECT 37.640 -13.890 37.810 -11.710 ;
        RECT 38.080 -12.660 38.250 -11.710 ;
        RECT 38.080 -12.830 38.290 -12.660 ;
        RECT 38.080 -13.710 38.250 -12.830 ;
        RECT 39.100 -13.890 39.270 -11.710 ;
        RECT 39.540 -12.660 39.710 -11.710 ;
        RECT 40.070 -12.660 40.240 -11.710 ;
        RECT 39.540 -12.830 40.240 -12.660 ;
        RECT 39.540 -13.710 39.710 -12.830 ;
        RECT 40.070 -13.710 40.240 -12.830 ;
        RECT 37.640 -14.060 39.270 -13.890 ;
        RECT 40.510 -13.890 40.680 -11.710 ;
        RECT 41.500 -12.660 41.670 -11.710 ;
        RECT 41.460 -12.830 41.670 -12.660 ;
        RECT 41.500 -13.710 41.670 -12.830 ;
        RECT 41.940 -13.890 42.110 -11.710 ;
        RECT 40.510 -13.950 42.110 -13.890 ;
        RECT 33.700 -14.120 34.930 -14.060 ;
        RECT 29.580 -14.490 29.910 -14.320 ;
        RECT 30.120 -14.490 30.450 -14.320 ;
        RECT 32.080 -14.490 32.410 -14.320 ;
        RECT 32.620 -14.490 32.950 -14.320 ;
        RECT 33.350 -14.460 34.590 -14.290 ;
        RECT 29.530 -17.700 29.700 -14.700 ;
        RECT 29.970 -18.180 30.140 -14.700 ;
        RECT 26.640 -18.350 30.140 -18.180 ;
        RECT 32.390 -18.180 32.560 -14.700 ;
        RECT 32.830 -17.700 33.000 -14.700 ;
        RECT 33.350 -17.700 33.520 -14.460 ;
        RECT 33.790 -17.700 33.960 -14.700 ;
        RECT 34.320 -17.700 34.490 -14.700 ;
        RECT 34.760 -17.700 34.930 -14.120 ;
        RECT 39.100 -14.290 39.270 -14.060 ;
        RECT 39.450 -14.060 42.110 -13.950 ;
        RECT 43.390 -13.890 43.560 -11.710 ;
        RECT 43.830 -12.660 44.000 -11.710 ;
        RECT 43.830 -12.830 44.040 -12.660 ;
        RECT 43.830 -13.710 44.000 -12.830 ;
        RECT 44.850 -13.890 45.020 -11.710 ;
        RECT 45.290 -12.660 45.460 -11.710 ;
        RECT 45.820 -12.660 45.990 -11.710 ;
        RECT 45.290 -12.830 45.990 -12.660 ;
        RECT 45.290 -13.710 45.460 -12.830 ;
        RECT 45.820 -13.710 45.990 -12.830 ;
        RECT 43.390 -14.060 45.020 -13.890 ;
        RECT 46.260 -13.890 46.430 -11.710 ;
        RECT 47.250 -12.660 47.420 -11.710 ;
        RECT 47.210 -12.830 47.420 -12.660 ;
        RECT 47.250 -13.710 47.420 -12.830 ;
        RECT 47.690 -13.890 47.860 -11.710 ;
        RECT 46.260 -13.950 47.860 -13.890 ;
        RECT 39.450 -14.120 40.680 -14.060 ;
        RECT 35.330 -14.490 35.660 -14.320 ;
        RECT 35.870 -14.490 36.200 -14.320 ;
        RECT 37.830 -14.490 38.160 -14.320 ;
        RECT 38.370 -14.490 38.700 -14.320 ;
        RECT 39.100 -14.460 40.340 -14.290 ;
        RECT 35.280 -17.700 35.450 -14.700 ;
        RECT 35.720 -18.180 35.890 -14.700 ;
        RECT 32.390 -18.350 35.890 -18.180 ;
        RECT 38.140 -18.180 38.310 -14.700 ;
        RECT 38.580 -17.700 38.750 -14.700 ;
        RECT 39.100 -17.700 39.270 -14.460 ;
        RECT 39.540 -17.700 39.710 -14.700 ;
        RECT 40.070 -17.700 40.240 -14.700 ;
        RECT 40.510 -17.700 40.680 -14.120 ;
        RECT 44.850 -14.290 45.020 -14.060 ;
        RECT 45.200 -14.060 47.860 -13.950 ;
        RECT 49.140 -13.890 49.310 -11.710 ;
        RECT 49.580 -12.660 49.750 -11.710 ;
        RECT 49.580 -12.830 49.790 -12.660 ;
        RECT 49.580 -13.710 49.750 -12.830 ;
        RECT 50.600 -13.890 50.770 -11.710 ;
        RECT 51.040 -12.660 51.210 -11.710 ;
        RECT 51.570 -12.660 51.740 -11.710 ;
        RECT 51.040 -12.830 51.740 -12.660 ;
        RECT 51.040 -13.710 51.210 -12.830 ;
        RECT 51.570 -13.710 51.740 -12.830 ;
        RECT 49.140 -14.060 50.770 -13.890 ;
        RECT 52.010 -13.890 52.180 -11.710 ;
        RECT 53.000 -12.660 53.170 -11.710 ;
        RECT 52.960 -12.830 53.170 -12.660 ;
        RECT 53.000 -13.710 53.170 -12.830 ;
        RECT 53.440 -13.890 53.610 -11.710 ;
        RECT 52.010 -13.950 53.610 -13.890 ;
        RECT 45.200 -14.120 46.430 -14.060 ;
        RECT 41.080 -14.490 41.410 -14.320 ;
        RECT 41.620 -14.490 41.950 -14.320 ;
        RECT 43.580 -14.490 43.910 -14.320 ;
        RECT 44.120 -14.490 44.450 -14.320 ;
        RECT 44.850 -14.460 46.090 -14.290 ;
        RECT 41.030 -17.700 41.200 -14.700 ;
        RECT 41.470 -18.180 41.640 -14.700 ;
        RECT 38.140 -18.350 41.640 -18.180 ;
        RECT 43.890 -18.180 44.060 -14.700 ;
        RECT 44.330 -17.700 44.500 -14.700 ;
        RECT 44.850 -17.700 45.020 -14.460 ;
        RECT 45.290 -17.700 45.460 -14.700 ;
        RECT 45.820 -17.700 45.990 -14.700 ;
        RECT 46.260 -17.700 46.430 -14.120 ;
        RECT 50.600 -14.290 50.770 -14.060 ;
        RECT 50.950 -14.060 53.610 -13.950 ;
        RECT 54.890 -13.890 55.060 -11.710 ;
        RECT 55.330 -12.660 55.500 -11.710 ;
        RECT 55.330 -12.830 55.540 -12.660 ;
        RECT 55.330 -13.710 55.500 -12.830 ;
        RECT 56.350 -13.890 56.520 -11.710 ;
        RECT 56.790 -12.660 56.960 -11.710 ;
        RECT 57.320 -12.660 57.490 -11.710 ;
        RECT 56.790 -12.830 57.490 -12.660 ;
        RECT 56.790 -13.710 56.960 -12.830 ;
        RECT 57.320 -13.710 57.490 -12.830 ;
        RECT 54.890 -14.060 56.520 -13.890 ;
        RECT 57.760 -13.890 57.930 -11.710 ;
        RECT 58.750 -12.660 58.920 -11.710 ;
        RECT 58.710 -12.830 58.920 -12.660 ;
        RECT 58.750 -13.710 58.920 -12.830 ;
        RECT 59.190 -13.890 59.360 -11.710 ;
        RECT 57.760 -13.950 59.360 -13.890 ;
        RECT 50.950 -14.120 52.180 -14.060 ;
        RECT 46.830 -14.490 47.160 -14.320 ;
        RECT 47.370 -14.490 47.700 -14.320 ;
        RECT 49.330 -14.490 49.660 -14.320 ;
        RECT 49.870 -14.490 50.200 -14.320 ;
        RECT 50.600 -14.460 51.840 -14.290 ;
        RECT 46.780 -17.700 46.950 -14.700 ;
        RECT 47.220 -18.180 47.390 -14.700 ;
        RECT 43.890 -18.350 47.390 -18.180 ;
        RECT 49.640 -18.180 49.810 -14.700 ;
        RECT 50.080 -17.700 50.250 -14.700 ;
        RECT 50.600 -17.700 50.770 -14.460 ;
        RECT 51.040 -17.700 51.210 -14.700 ;
        RECT 51.570 -17.700 51.740 -14.700 ;
        RECT 52.010 -17.700 52.180 -14.120 ;
        RECT 56.350 -14.290 56.520 -14.060 ;
        RECT 56.700 -14.060 59.360 -13.950 ;
        RECT 60.640 -13.890 60.810 -11.710 ;
        RECT 61.080 -12.660 61.250 -11.710 ;
        RECT 61.080 -12.830 61.290 -12.660 ;
        RECT 61.080 -13.710 61.250 -12.830 ;
        RECT 62.100 -13.890 62.270 -11.710 ;
        RECT 62.540 -12.660 62.710 -11.710 ;
        RECT 63.070 -12.660 63.240 -11.710 ;
        RECT 62.540 -12.830 63.240 -12.660 ;
        RECT 62.540 -13.710 62.710 -12.830 ;
        RECT 63.070 -13.710 63.240 -12.830 ;
        RECT 60.640 -14.060 62.270 -13.890 ;
        RECT 63.510 -13.890 63.680 -11.710 ;
        RECT 64.500 -12.660 64.670 -11.710 ;
        RECT 64.460 -12.830 64.670 -12.660 ;
        RECT 64.500 -13.710 64.670 -12.830 ;
        RECT 64.940 -13.890 65.110 -11.710 ;
        RECT 63.510 -13.950 65.110 -13.890 ;
        RECT 56.700 -14.120 57.930 -14.060 ;
        RECT 52.580 -14.490 52.910 -14.320 ;
        RECT 53.120 -14.490 53.450 -14.320 ;
        RECT 55.080 -14.490 55.410 -14.320 ;
        RECT 55.620 -14.490 55.950 -14.320 ;
        RECT 56.350 -14.460 57.590 -14.290 ;
        RECT 52.530 -17.700 52.700 -14.700 ;
        RECT 52.970 -18.180 53.140 -14.700 ;
        RECT 49.640 -18.350 53.140 -18.180 ;
        RECT 55.390 -18.180 55.560 -14.700 ;
        RECT 55.830 -17.700 56.000 -14.700 ;
        RECT 56.350 -17.700 56.520 -14.460 ;
        RECT 56.790 -17.700 56.960 -14.700 ;
        RECT 57.320 -17.700 57.490 -14.700 ;
        RECT 57.760 -17.700 57.930 -14.120 ;
        RECT 62.100 -14.290 62.270 -14.060 ;
        RECT 62.450 -14.060 65.110 -13.950 ;
        RECT 66.390 -13.890 66.560 -11.710 ;
        RECT 66.830 -12.660 67.000 -11.710 ;
        RECT 66.830 -12.830 67.040 -12.660 ;
        RECT 66.830 -13.710 67.000 -12.830 ;
        RECT 67.850 -13.890 68.020 -11.710 ;
        RECT 68.290 -12.660 68.460 -11.710 ;
        RECT 68.820 -12.660 68.990 -11.710 ;
        RECT 68.290 -12.830 68.990 -12.660 ;
        RECT 68.290 -13.710 68.460 -12.830 ;
        RECT 68.820 -13.710 68.990 -12.830 ;
        RECT 66.390 -14.060 68.020 -13.890 ;
        RECT 69.260 -13.890 69.430 -11.710 ;
        RECT 70.250 -12.660 70.420 -11.710 ;
        RECT 70.210 -12.830 70.420 -12.660 ;
        RECT 70.250 -13.710 70.420 -12.830 ;
        RECT 70.690 -13.890 70.860 -11.710 ;
        RECT 69.260 -13.950 70.860 -13.890 ;
        RECT 62.450 -14.120 63.680 -14.060 ;
        RECT 58.330 -14.490 58.660 -14.320 ;
        RECT 58.870 -14.490 59.200 -14.320 ;
        RECT 60.830 -14.490 61.160 -14.320 ;
        RECT 61.370 -14.490 61.700 -14.320 ;
        RECT 62.100 -14.460 63.340 -14.290 ;
        RECT 58.280 -17.700 58.450 -14.700 ;
        RECT 58.720 -18.180 58.890 -14.700 ;
        RECT 55.390 -18.350 58.890 -18.180 ;
        RECT 61.140 -18.180 61.310 -14.700 ;
        RECT 61.580 -17.700 61.750 -14.700 ;
        RECT 62.100 -17.700 62.270 -14.460 ;
        RECT 62.540 -17.700 62.710 -14.700 ;
        RECT 63.070 -17.700 63.240 -14.700 ;
        RECT 63.510 -17.700 63.680 -14.120 ;
        RECT 67.850 -14.290 68.020 -14.060 ;
        RECT 68.200 -14.060 70.860 -13.950 ;
        RECT 72.140 -13.890 72.310 -11.710 ;
        RECT 72.580 -12.660 72.750 -11.710 ;
        RECT 72.580 -12.830 72.790 -12.660 ;
        RECT 72.580 -13.710 72.750 -12.830 ;
        RECT 73.600 -13.890 73.770 -11.710 ;
        RECT 74.040 -12.660 74.210 -11.710 ;
        RECT 74.570 -12.660 74.740 -11.710 ;
        RECT 74.040 -12.830 74.740 -12.660 ;
        RECT 74.040 -13.710 74.210 -12.830 ;
        RECT 74.570 -13.710 74.740 -12.830 ;
        RECT 72.140 -14.060 73.770 -13.890 ;
        RECT 75.010 -13.890 75.180 -11.710 ;
        RECT 76.000 -12.660 76.170 -11.710 ;
        RECT 75.960 -12.830 76.170 -12.660 ;
        RECT 76.000 -13.710 76.170 -12.830 ;
        RECT 76.440 -13.890 76.610 -11.710 ;
        RECT 75.010 -13.950 76.610 -13.890 ;
        RECT 68.200 -14.120 69.430 -14.060 ;
        RECT 64.080 -14.490 64.410 -14.320 ;
        RECT 64.620 -14.490 64.950 -14.320 ;
        RECT 66.580 -14.490 66.910 -14.320 ;
        RECT 67.120 -14.490 67.450 -14.320 ;
        RECT 67.850 -14.460 69.090 -14.290 ;
        RECT 64.030 -17.700 64.200 -14.700 ;
        RECT 64.470 -18.180 64.640 -14.700 ;
        RECT 61.140 -18.350 64.640 -18.180 ;
        RECT 66.890 -18.180 67.060 -14.700 ;
        RECT 67.330 -17.700 67.500 -14.700 ;
        RECT 67.850 -17.700 68.020 -14.460 ;
        RECT 68.290 -17.700 68.460 -14.700 ;
        RECT 68.820 -17.700 68.990 -14.700 ;
        RECT 69.260 -17.700 69.430 -14.120 ;
        RECT 73.600 -14.290 73.770 -14.060 ;
        RECT 73.950 -14.060 76.610 -13.950 ;
        RECT 77.890 -13.890 78.060 -11.710 ;
        RECT 78.330 -12.660 78.500 -11.710 ;
        RECT 78.330 -12.830 78.540 -12.660 ;
        RECT 78.330 -13.710 78.500 -12.830 ;
        RECT 79.350 -13.890 79.520 -11.710 ;
        RECT 79.790 -12.660 79.960 -11.710 ;
        RECT 80.320 -12.660 80.490 -11.710 ;
        RECT 79.790 -12.830 80.490 -12.660 ;
        RECT 79.790 -13.710 79.960 -12.830 ;
        RECT 80.320 -13.710 80.490 -12.830 ;
        RECT 77.890 -14.060 79.520 -13.890 ;
        RECT 80.760 -13.890 80.930 -11.710 ;
        RECT 81.750 -12.660 81.920 -11.710 ;
        RECT 81.710 -12.830 81.920 -12.660 ;
        RECT 81.750 -13.710 81.920 -12.830 ;
        RECT 82.190 -13.890 82.360 -11.710 ;
        RECT 80.760 -13.950 82.360 -13.890 ;
        RECT 73.950 -14.120 75.180 -14.060 ;
        RECT 69.830 -14.490 70.160 -14.320 ;
        RECT 70.370 -14.490 70.700 -14.320 ;
        RECT 72.330 -14.490 72.660 -14.320 ;
        RECT 72.870 -14.490 73.200 -14.320 ;
        RECT 73.600 -14.460 74.840 -14.290 ;
        RECT 69.780 -17.700 69.950 -14.700 ;
        RECT 70.220 -18.180 70.390 -14.700 ;
        RECT 66.890 -18.350 70.390 -18.180 ;
        RECT 72.640 -18.180 72.810 -14.700 ;
        RECT 73.080 -17.700 73.250 -14.700 ;
        RECT 73.600 -17.700 73.770 -14.460 ;
        RECT 74.040 -17.700 74.210 -14.700 ;
        RECT 74.570 -17.700 74.740 -14.700 ;
        RECT 75.010 -17.700 75.180 -14.120 ;
        RECT 79.350 -14.290 79.520 -14.060 ;
        RECT 79.700 -14.060 82.360 -13.950 ;
        RECT 83.640 -13.890 83.810 -11.710 ;
        RECT 84.080 -12.660 84.250 -11.710 ;
        RECT 84.080 -12.830 84.290 -12.660 ;
        RECT 84.080 -13.710 84.250 -12.830 ;
        RECT 85.100 -13.890 85.270 -11.710 ;
        RECT 85.540 -12.660 85.710 -11.710 ;
        RECT 86.070 -12.660 86.240 -11.710 ;
        RECT 85.540 -12.830 86.240 -12.660 ;
        RECT 85.540 -13.710 85.710 -12.830 ;
        RECT 86.070 -13.710 86.240 -12.830 ;
        RECT 83.640 -14.060 85.270 -13.890 ;
        RECT 86.510 -13.890 86.680 -11.710 ;
        RECT 87.500 -12.660 87.670 -11.710 ;
        RECT 87.460 -12.830 87.670 -12.660 ;
        RECT 87.500 -13.710 87.670 -12.830 ;
        RECT 87.940 -13.890 88.110 -11.710 ;
        RECT 86.510 -13.950 88.110 -13.890 ;
        RECT 79.700 -14.120 80.930 -14.060 ;
        RECT 75.580 -14.490 75.910 -14.320 ;
        RECT 76.120 -14.490 76.450 -14.320 ;
        RECT 78.080 -14.490 78.410 -14.320 ;
        RECT 78.620 -14.490 78.950 -14.320 ;
        RECT 79.350 -14.460 80.590 -14.290 ;
        RECT 75.530 -17.700 75.700 -14.700 ;
        RECT 75.970 -18.180 76.140 -14.700 ;
        RECT 72.640 -18.350 76.140 -18.180 ;
        RECT 78.390 -18.180 78.560 -14.700 ;
        RECT 78.830 -17.700 79.000 -14.700 ;
        RECT 79.350 -17.700 79.520 -14.460 ;
        RECT 79.790 -17.700 79.960 -14.700 ;
        RECT 80.320 -17.700 80.490 -14.700 ;
        RECT 80.760 -17.700 80.930 -14.120 ;
        RECT 85.100 -14.290 85.270 -14.060 ;
        RECT 85.450 -14.060 88.110 -13.950 ;
        RECT 89.390 -13.890 89.560 -11.710 ;
        RECT 89.830 -12.660 90.000 -11.710 ;
        RECT 89.830 -12.830 90.040 -12.660 ;
        RECT 89.830 -13.710 90.000 -12.830 ;
        RECT 90.850 -13.890 91.020 -11.710 ;
        RECT 91.290 -12.660 91.460 -11.710 ;
        RECT 91.820 -12.660 91.990 -11.710 ;
        RECT 91.290 -12.830 91.990 -12.660 ;
        RECT 91.290 -13.710 91.460 -12.830 ;
        RECT 91.820 -13.710 91.990 -12.830 ;
        RECT 89.390 -14.060 91.020 -13.890 ;
        RECT 92.260 -13.890 92.430 -11.710 ;
        RECT 93.250 -12.660 93.420 -11.710 ;
        RECT 93.210 -12.830 93.420 -12.660 ;
        RECT 93.250 -13.710 93.420 -12.830 ;
        RECT 93.690 -13.890 93.860 -11.710 ;
        RECT 92.260 -13.950 93.860 -13.890 ;
        RECT 85.450 -14.120 86.680 -14.060 ;
        RECT 81.330 -14.490 81.660 -14.320 ;
        RECT 81.870 -14.490 82.200 -14.320 ;
        RECT 83.830 -14.490 84.160 -14.320 ;
        RECT 84.370 -14.490 84.700 -14.320 ;
        RECT 85.100 -14.460 86.340 -14.290 ;
        RECT 81.280 -17.700 81.450 -14.700 ;
        RECT 81.720 -18.180 81.890 -14.700 ;
        RECT 78.390 -18.350 81.890 -18.180 ;
        RECT 84.140 -18.180 84.310 -14.700 ;
        RECT 84.580 -17.700 84.750 -14.700 ;
        RECT 85.100 -17.700 85.270 -14.460 ;
        RECT 85.540 -17.700 85.710 -14.700 ;
        RECT 86.070 -17.700 86.240 -14.700 ;
        RECT 86.510 -17.700 86.680 -14.120 ;
        RECT 90.850 -14.290 91.020 -14.060 ;
        RECT 91.200 -14.060 93.860 -13.950 ;
        RECT 91.200 -14.120 92.430 -14.060 ;
        RECT 87.080 -14.490 87.410 -14.320 ;
        RECT 87.620 -14.490 87.950 -14.320 ;
        RECT 89.580 -14.490 89.910 -14.320 ;
        RECT 90.120 -14.490 90.450 -14.320 ;
        RECT 90.850 -14.460 92.090 -14.290 ;
        RECT 87.030 -17.700 87.200 -14.700 ;
        RECT 87.470 -18.180 87.640 -14.700 ;
        RECT 84.140 -18.350 87.640 -18.180 ;
        RECT 89.890 -18.180 90.060 -14.700 ;
        RECT 90.330 -17.700 90.500 -14.700 ;
        RECT 90.850 -17.700 91.020 -14.460 ;
        RECT 91.290 -17.700 91.460 -14.700 ;
        RECT 91.820 -17.700 91.990 -14.700 ;
        RECT 92.260 -17.700 92.430 -14.120 ;
        RECT 92.830 -14.490 93.160 -14.320 ;
        RECT 93.370 -14.490 93.700 -14.320 ;
        RECT 92.780 -17.700 92.950 -14.700 ;
        RECT 93.220 -18.180 93.390 -14.700 ;
        RECT 89.890 -18.350 93.390 -18.180 ;
        RECT 3.400 -18.690 3.730 -18.520 ;
        RECT 3.900 -18.790 6.900 -18.620 ;
        RECT 7.080 -18.700 7.410 -18.530 ;
        RECT 9.150 -18.690 9.480 -18.520 ;
        RECT 9.650 -18.790 12.650 -18.620 ;
        RECT 12.830 -18.700 13.160 -18.530 ;
        RECT 14.900 -18.690 15.230 -18.520 ;
        RECT 15.400 -18.790 18.400 -18.620 ;
        RECT 18.580 -18.700 18.910 -18.530 ;
        RECT 20.650 -18.690 20.980 -18.520 ;
        RECT 21.150 -18.790 24.150 -18.620 ;
        RECT 24.330 -18.700 24.660 -18.530 ;
        RECT 26.400 -18.690 26.730 -18.520 ;
        RECT 26.900 -18.790 29.900 -18.620 ;
        RECT 30.080 -18.700 30.410 -18.530 ;
        RECT 32.150 -18.690 32.480 -18.520 ;
        RECT 32.650 -18.790 35.650 -18.620 ;
        RECT 35.830 -18.700 36.160 -18.530 ;
        RECT 37.900 -18.690 38.230 -18.520 ;
        RECT 38.400 -18.790 41.400 -18.620 ;
        RECT 41.580 -18.700 41.910 -18.530 ;
        RECT 43.650 -18.690 43.980 -18.520 ;
        RECT 44.150 -18.790 47.150 -18.620 ;
        RECT 47.330 -18.700 47.660 -18.530 ;
        RECT 49.400 -18.690 49.730 -18.520 ;
        RECT 49.900 -18.790 52.900 -18.620 ;
        RECT 53.080 -18.700 53.410 -18.530 ;
        RECT 55.150 -18.690 55.480 -18.520 ;
        RECT 55.650 -18.790 58.650 -18.620 ;
        RECT 58.830 -18.700 59.160 -18.530 ;
        RECT 60.900 -18.690 61.230 -18.520 ;
        RECT 61.400 -18.790 64.400 -18.620 ;
        RECT 64.580 -18.700 64.910 -18.530 ;
        RECT 66.650 -18.690 66.980 -18.520 ;
        RECT 67.150 -18.790 70.150 -18.620 ;
        RECT 70.330 -18.700 70.660 -18.530 ;
        RECT 72.400 -18.690 72.730 -18.520 ;
        RECT 72.900 -18.790 75.900 -18.620 ;
        RECT 76.080 -18.700 76.410 -18.530 ;
        RECT 78.150 -18.690 78.480 -18.520 ;
        RECT 78.650 -18.790 81.650 -18.620 ;
        RECT 81.830 -18.700 82.160 -18.530 ;
        RECT 83.900 -18.690 84.230 -18.520 ;
        RECT 84.400 -18.790 87.400 -18.620 ;
        RECT 87.580 -18.700 87.910 -18.530 ;
        RECT 89.650 -18.690 89.980 -18.520 ;
        RECT 90.150 -18.790 93.150 -18.620 ;
        RECT 93.330 -18.700 93.660 -18.530 ;
        RECT 5.390 -19.130 5.560 -18.790 ;
        RECT 8.000 -19.130 8.410 -18.960 ;
        RECT 11.140 -19.130 11.310 -18.790 ;
        RECT 13.750 -19.130 14.160 -18.960 ;
        RECT 16.890 -19.130 17.060 -18.790 ;
        RECT 19.500 -19.130 19.910 -18.960 ;
        RECT 22.640 -19.130 22.810 -18.790 ;
        RECT 25.250 -19.130 25.660 -18.960 ;
        RECT 28.390 -19.130 28.560 -18.790 ;
        RECT 31.000 -19.130 31.410 -18.960 ;
        RECT 34.140 -19.130 34.310 -18.790 ;
        RECT 36.750 -19.130 37.160 -18.960 ;
        RECT 39.890 -19.130 40.060 -18.790 ;
        RECT 42.500 -19.130 42.910 -18.960 ;
        RECT 45.640 -19.130 45.810 -18.790 ;
        RECT 48.250 -19.130 48.660 -18.960 ;
        RECT 51.390 -19.130 51.560 -18.790 ;
        RECT 54.000 -19.130 54.410 -18.960 ;
        RECT 57.140 -19.130 57.310 -18.790 ;
        RECT 59.750 -19.130 60.160 -18.960 ;
        RECT 62.890 -19.130 63.060 -18.790 ;
        RECT 65.500 -19.130 65.910 -18.960 ;
        RECT 68.640 -19.130 68.810 -18.790 ;
        RECT 71.250 -19.130 71.660 -18.960 ;
        RECT 74.390 -19.130 74.560 -18.790 ;
        RECT 77.000 -19.130 77.410 -18.960 ;
        RECT 80.140 -19.130 80.310 -18.790 ;
        RECT 82.750 -19.130 83.160 -18.960 ;
        RECT 85.890 -19.130 86.060 -18.790 ;
        RECT 88.500 -19.130 88.910 -18.960 ;
        RECT 91.640 -19.130 91.810 -18.790 ;
        RECT 94.110 -19.130 94.520 -18.960 ;
        RECT 4.350 -19.480 4.520 -19.440 ;
        RECT 6.230 -19.480 6.400 -19.440 ;
        RECT 10.100 -19.480 10.270 -19.440 ;
        RECT 11.980 -19.480 12.150 -19.440 ;
        RECT 15.850 -19.480 16.020 -19.440 ;
        RECT 17.730 -19.480 17.900 -19.440 ;
        RECT 21.600 -19.480 21.770 -19.440 ;
        RECT 23.480 -19.480 23.650 -19.440 ;
        RECT 27.350 -19.480 27.520 -19.440 ;
        RECT 29.230 -19.480 29.400 -19.440 ;
        RECT 33.100 -19.480 33.270 -19.440 ;
        RECT 34.980 -19.480 35.150 -19.440 ;
        RECT 38.850 -19.480 39.020 -19.440 ;
        RECT 40.730 -19.480 40.900 -19.440 ;
        RECT 44.600 -19.480 44.770 -19.440 ;
        RECT 46.480 -19.480 46.650 -19.440 ;
        RECT 50.350 -19.480 50.520 -19.440 ;
        RECT 52.230 -19.480 52.400 -19.440 ;
        RECT 56.100 -19.480 56.270 -19.440 ;
        RECT 57.980 -19.480 58.150 -19.440 ;
        RECT 61.850 -19.480 62.020 -19.440 ;
        RECT 63.730 -19.480 63.900 -19.440 ;
        RECT 67.600 -19.480 67.770 -19.440 ;
        RECT 69.480 -19.480 69.650 -19.440 ;
        RECT 73.350 -19.480 73.520 -19.440 ;
        RECT 75.230 -19.480 75.400 -19.440 ;
        RECT 79.100 -19.480 79.270 -19.440 ;
        RECT 80.980 -19.480 81.150 -19.440 ;
        RECT 84.850 -19.480 85.020 -19.440 ;
        RECT 86.730 -19.480 86.900 -19.440 ;
        RECT 90.600 -19.480 90.770 -19.440 ;
        RECT 92.480 -19.480 92.650 -19.440 ;
        RECT 4.270 -19.650 4.600 -19.480 ;
        RECT 6.150 -19.650 6.480 -19.480 ;
        RECT 10.020 -19.650 10.350 -19.480 ;
        RECT 11.900 -19.650 12.230 -19.480 ;
        RECT 15.770 -19.650 16.100 -19.480 ;
        RECT 17.650 -19.650 17.980 -19.480 ;
        RECT 21.520 -19.650 21.850 -19.480 ;
        RECT 23.400 -19.650 23.730 -19.480 ;
        RECT 27.270 -19.650 27.600 -19.480 ;
        RECT 29.150 -19.650 29.480 -19.480 ;
        RECT 33.020 -19.650 33.350 -19.480 ;
        RECT 34.900 -19.650 35.230 -19.480 ;
        RECT 38.770 -19.650 39.100 -19.480 ;
        RECT 40.650 -19.650 40.980 -19.480 ;
        RECT 44.520 -19.650 44.850 -19.480 ;
        RECT 46.400 -19.650 46.730 -19.480 ;
        RECT 50.270 -19.650 50.600 -19.480 ;
        RECT 52.150 -19.650 52.480 -19.480 ;
        RECT 56.020 -19.650 56.350 -19.480 ;
        RECT 57.900 -19.650 58.230 -19.480 ;
        RECT 61.770 -19.650 62.100 -19.480 ;
        RECT 63.650 -19.650 63.980 -19.480 ;
        RECT 67.520 -19.650 67.850 -19.480 ;
        RECT 69.400 -19.650 69.730 -19.480 ;
        RECT 73.270 -19.650 73.600 -19.480 ;
        RECT 75.150 -19.650 75.480 -19.480 ;
        RECT 79.020 -19.650 79.350 -19.480 ;
        RECT 80.900 -19.650 81.230 -19.480 ;
        RECT 84.770 -19.650 85.100 -19.480 ;
        RECT 86.650 -19.650 86.980 -19.480 ;
        RECT 90.520 -19.650 90.850 -19.480 ;
        RECT 92.400 -19.650 92.730 -19.480 ;
        RECT 4.350 -19.690 4.520 -19.650 ;
        RECT 6.230 -19.690 6.400 -19.650 ;
        RECT 10.100 -19.690 10.270 -19.650 ;
        RECT 11.980 -19.690 12.150 -19.650 ;
        RECT 15.850 -19.690 16.020 -19.650 ;
        RECT 17.730 -19.690 17.900 -19.650 ;
        RECT 21.600 -19.690 21.770 -19.650 ;
        RECT 23.480 -19.690 23.650 -19.650 ;
        RECT 27.350 -19.690 27.520 -19.650 ;
        RECT 29.230 -19.690 29.400 -19.650 ;
        RECT 33.100 -19.690 33.270 -19.650 ;
        RECT 34.980 -19.690 35.150 -19.650 ;
        RECT 38.850 -19.690 39.020 -19.650 ;
        RECT 40.730 -19.690 40.900 -19.650 ;
        RECT 44.600 -19.690 44.770 -19.650 ;
        RECT 46.480 -19.690 46.650 -19.650 ;
        RECT 50.350 -19.690 50.520 -19.650 ;
        RECT 52.230 -19.690 52.400 -19.650 ;
        RECT 56.100 -19.690 56.270 -19.650 ;
        RECT 57.980 -19.690 58.150 -19.650 ;
        RECT 61.850 -19.690 62.020 -19.650 ;
        RECT 63.730 -19.690 63.900 -19.650 ;
        RECT 67.600 -19.690 67.770 -19.650 ;
        RECT 69.480 -19.690 69.650 -19.650 ;
        RECT 73.350 -19.690 73.520 -19.650 ;
        RECT 75.230 -19.690 75.400 -19.650 ;
        RECT 79.100 -19.690 79.270 -19.650 ;
        RECT 80.980 -19.690 81.150 -19.650 ;
        RECT 84.850 -19.690 85.020 -19.650 ;
        RECT 86.730 -19.690 86.900 -19.650 ;
        RECT 90.600 -19.690 90.770 -19.650 ;
        RECT 92.480 -19.690 92.650 -19.650 ;
        RECT 3.140 -20.360 3.310 -20.230 ;
        RECT 3.100 -20.530 3.370 -20.360 ;
        RECT 3.140 -20.650 3.310 -20.530 ;
        RECT 3.120 -21.050 3.290 -21.010 ;
        RECT 3.580 -21.030 3.750 -20.230 ;
        RECT 4.150 -20.860 4.320 -19.860 ;
        RECT 4.590 -20.860 4.760 -19.860 ;
        RECT 5.030 -20.370 5.200 -19.860 ;
        RECT 5.550 -20.370 5.720 -19.860 ;
        RECT 4.970 -20.540 5.240 -20.370 ;
        RECT 5.510 -20.540 5.780 -20.370 ;
        RECT 5.030 -20.860 5.200 -20.540 ;
        RECT 5.550 -20.860 5.720 -20.540 ;
        RECT 5.990 -20.860 6.160 -19.860 ;
        RECT 6.430 -20.860 6.600 -19.860 ;
        RECT 3.040 -21.220 3.370 -21.050 ;
        RECT 3.580 -21.070 3.810 -21.030 ;
        RECT 3.120 -21.260 3.290 -21.220 ;
        RECT 3.580 -21.240 3.870 -21.070 ;
        RECT 4.750 -21.240 5.080 -21.070 ;
        RECT 5.670 -21.240 6.000 -21.070 ;
        RECT 3.580 -21.280 3.810 -21.240 ;
        RECT 3.140 -21.840 3.310 -21.500 ;
        RECT 3.100 -22.010 3.370 -21.840 ;
        RECT 3.140 -22.340 3.310 -22.010 ;
        RECT 3.580 -22.340 3.750 -21.280 ;
        RECT 4.830 -21.500 5.000 -21.240 ;
        RECT 7.000 -21.500 7.170 -20.230 ;
        RECT 7.440 -20.360 7.610 -20.230 ;
        RECT 8.890 -20.360 9.060 -20.230 ;
        RECT 7.380 -20.530 7.650 -20.360 ;
        RECT 8.850 -20.530 9.120 -20.360 ;
        RECT 7.440 -20.650 7.610 -20.530 ;
        RECT 8.890 -20.650 9.060 -20.530 ;
        RECT 7.450 -21.070 7.620 -21.030 ;
        RECT 8.870 -21.050 9.040 -21.010 ;
        RECT 9.330 -21.030 9.500 -20.230 ;
        RECT 9.900 -20.860 10.070 -19.860 ;
        RECT 10.340 -20.860 10.510 -19.860 ;
        RECT 10.780 -20.370 10.950 -19.860 ;
        RECT 11.300 -20.370 11.470 -19.860 ;
        RECT 10.720 -20.540 10.990 -20.370 ;
        RECT 11.260 -20.540 11.530 -20.370 ;
        RECT 10.780 -20.860 10.950 -20.540 ;
        RECT 11.300 -20.860 11.470 -20.540 ;
        RECT 11.740 -20.860 11.910 -19.860 ;
        RECT 12.180 -20.860 12.350 -19.860 ;
        RECT 7.370 -21.240 7.700 -21.070 ;
        RECT 8.790 -21.220 9.120 -21.050 ;
        RECT 9.330 -21.070 9.560 -21.030 ;
        RECT 7.450 -21.280 7.620 -21.240 ;
        RECT 8.870 -21.260 9.040 -21.220 ;
        RECT 9.330 -21.240 9.620 -21.070 ;
        RECT 10.500 -21.240 10.830 -21.070 ;
        RECT 11.420 -21.240 11.750 -21.070 ;
        RECT 9.330 -21.280 9.560 -21.240 ;
        RECT 4.830 -21.670 7.170 -21.500 ;
        RECT 7.000 -22.340 7.170 -21.670 ;
        RECT 7.440 -21.780 7.610 -21.500 ;
        RECT 7.420 -21.830 7.610 -21.780 ;
        RECT 7.420 -21.840 8.410 -21.830 ;
        RECT 8.890 -21.840 9.060 -21.500 ;
        RECT 7.380 -22.000 8.410 -21.840 ;
        RECT 7.380 -22.010 7.650 -22.000 ;
        RECT 8.850 -22.010 9.120 -21.840 ;
        RECT 7.420 -22.070 7.610 -22.010 ;
        RECT 7.440 -22.340 7.610 -22.070 ;
        RECT 8.890 -22.340 9.060 -22.010 ;
        RECT 9.330 -22.340 9.500 -21.280 ;
        RECT 10.580 -21.500 10.750 -21.240 ;
        RECT 12.750 -21.500 12.920 -20.230 ;
        RECT 13.190 -20.360 13.360 -20.230 ;
        RECT 14.640 -20.360 14.810 -20.230 ;
        RECT 13.130 -20.530 13.400 -20.360 ;
        RECT 14.600 -20.530 14.870 -20.360 ;
        RECT 13.190 -20.650 13.360 -20.530 ;
        RECT 14.640 -20.650 14.810 -20.530 ;
        RECT 13.200 -21.070 13.370 -21.030 ;
        RECT 14.620 -21.050 14.790 -21.010 ;
        RECT 15.080 -21.030 15.250 -20.230 ;
        RECT 15.650 -20.860 15.820 -19.860 ;
        RECT 16.090 -20.860 16.260 -19.860 ;
        RECT 16.530 -20.370 16.700 -19.860 ;
        RECT 17.050 -20.370 17.220 -19.860 ;
        RECT 16.470 -20.540 16.740 -20.370 ;
        RECT 17.010 -20.540 17.280 -20.370 ;
        RECT 16.530 -20.860 16.700 -20.540 ;
        RECT 17.050 -20.860 17.220 -20.540 ;
        RECT 17.490 -20.860 17.660 -19.860 ;
        RECT 17.930 -20.860 18.100 -19.860 ;
        RECT 13.120 -21.240 13.450 -21.070 ;
        RECT 14.540 -21.220 14.870 -21.050 ;
        RECT 15.080 -21.070 15.310 -21.030 ;
        RECT 13.200 -21.280 13.370 -21.240 ;
        RECT 14.620 -21.260 14.790 -21.220 ;
        RECT 15.080 -21.240 15.370 -21.070 ;
        RECT 16.250 -21.240 16.580 -21.070 ;
        RECT 17.170 -21.240 17.500 -21.070 ;
        RECT 15.080 -21.280 15.310 -21.240 ;
        RECT 10.580 -21.670 12.920 -21.500 ;
        RECT 12.750 -22.340 12.920 -21.670 ;
        RECT 13.190 -21.780 13.360 -21.500 ;
        RECT 13.170 -21.840 13.360 -21.780 ;
        RECT 14.640 -21.840 14.810 -21.500 ;
        RECT 13.130 -22.010 14.160 -21.840 ;
        RECT 14.600 -22.010 14.870 -21.840 ;
        RECT 13.170 -22.070 13.360 -22.010 ;
        RECT 13.190 -22.340 13.360 -22.070 ;
        RECT 14.640 -22.340 14.810 -22.010 ;
        RECT 15.080 -22.340 15.250 -21.280 ;
        RECT 16.330 -21.500 16.500 -21.240 ;
        RECT 18.500 -21.500 18.670 -20.230 ;
        RECT 18.940 -20.360 19.110 -20.230 ;
        RECT 20.390 -20.360 20.560 -20.230 ;
        RECT 18.880 -20.530 19.150 -20.360 ;
        RECT 20.350 -20.530 20.620 -20.360 ;
        RECT 18.940 -20.650 19.110 -20.530 ;
        RECT 20.390 -20.650 20.560 -20.530 ;
        RECT 18.950 -21.070 19.120 -21.030 ;
        RECT 20.370 -21.050 20.540 -21.010 ;
        RECT 20.830 -21.030 21.000 -20.230 ;
        RECT 21.400 -20.860 21.570 -19.860 ;
        RECT 21.840 -20.860 22.010 -19.860 ;
        RECT 22.280 -20.370 22.450 -19.860 ;
        RECT 22.800 -20.370 22.970 -19.860 ;
        RECT 22.220 -20.540 22.490 -20.370 ;
        RECT 22.760 -20.540 23.030 -20.370 ;
        RECT 22.280 -20.860 22.450 -20.540 ;
        RECT 22.800 -20.860 22.970 -20.540 ;
        RECT 23.240 -20.860 23.410 -19.860 ;
        RECT 23.680 -20.860 23.850 -19.860 ;
        RECT 18.870 -21.240 19.200 -21.070 ;
        RECT 20.290 -21.220 20.620 -21.050 ;
        RECT 20.830 -21.070 21.060 -21.030 ;
        RECT 18.950 -21.280 19.120 -21.240 ;
        RECT 20.370 -21.260 20.540 -21.220 ;
        RECT 20.830 -21.240 21.120 -21.070 ;
        RECT 22.000 -21.240 22.330 -21.070 ;
        RECT 22.920 -21.240 23.250 -21.070 ;
        RECT 20.830 -21.280 21.060 -21.240 ;
        RECT 16.330 -21.670 18.670 -21.500 ;
        RECT 18.500 -22.340 18.670 -21.670 ;
        RECT 18.940 -21.780 19.110 -21.500 ;
        RECT 18.920 -21.840 19.110 -21.780 ;
        RECT 20.390 -21.840 20.560 -21.500 ;
        RECT 18.880 -22.010 19.910 -21.840 ;
        RECT 20.350 -22.010 20.620 -21.840 ;
        RECT 18.920 -22.070 19.110 -22.010 ;
        RECT 18.940 -22.340 19.110 -22.070 ;
        RECT 20.390 -22.340 20.560 -22.010 ;
        RECT 20.830 -22.340 21.000 -21.280 ;
        RECT 22.080 -21.500 22.250 -21.240 ;
        RECT 24.250 -21.500 24.420 -20.230 ;
        RECT 24.690 -20.360 24.860 -20.230 ;
        RECT 26.140 -20.360 26.310 -20.230 ;
        RECT 24.630 -20.530 24.900 -20.360 ;
        RECT 26.100 -20.530 26.370 -20.360 ;
        RECT 24.690 -20.650 24.860 -20.530 ;
        RECT 26.140 -20.650 26.310 -20.530 ;
        RECT 24.700 -21.070 24.870 -21.030 ;
        RECT 26.120 -21.050 26.290 -21.010 ;
        RECT 26.580 -21.030 26.750 -20.230 ;
        RECT 27.150 -20.860 27.320 -19.860 ;
        RECT 27.590 -20.860 27.760 -19.860 ;
        RECT 28.030 -20.370 28.200 -19.860 ;
        RECT 28.550 -20.370 28.720 -19.860 ;
        RECT 27.970 -20.540 28.240 -20.370 ;
        RECT 28.510 -20.540 28.780 -20.370 ;
        RECT 28.030 -20.860 28.200 -20.540 ;
        RECT 28.550 -20.860 28.720 -20.540 ;
        RECT 28.990 -20.860 29.160 -19.860 ;
        RECT 29.430 -20.860 29.600 -19.860 ;
        RECT 24.620 -21.240 24.950 -21.070 ;
        RECT 26.040 -21.220 26.370 -21.050 ;
        RECT 26.580 -21.070 26.810 -21.030 ;
        RECT 24.700 -21.280 24.870 -21.240 ;
        RECT 26.120 -21.260 26.290 -21.220 ;
        RECT 26.580 -21.240 26.870 -21.070 ;
        RECT 27.750 -21.240 28.080 -21.070 ;
        RECT 28.670 -21.240 29.000 -21.070 ;
        RECT 26.580 -21.280 26.810 -21.240 ;
        RECT 22.080 -21.670 24.420 -21.500 ;
        RECT 24.250 -22.340 24.420 -21.670 ;
        RECT 24.690 -21.780 24.860 -21.500 ;
        RECT 24.670 -21.840 24.860 -21.780 ;
        RECT 26.140 -21.840 26.310 -21.500 ;
        RECT 24.630 -22.010 25.660 -21.840 ;
        RECT 26.100 -22.010 26.370 -21.840 ;
        RECT 24.670 -22.070 24.860 -22.010 ;
        RECT 24.690 -22.340 24.860 -22.070 ;
        RECT 26.140 -22.340 26.310 -22.010 ;
        RECT 26.580 -22.340 26.750 -21.280 ;
        RECT 27.830 -21.500 28.000 -21.240 ;
        RECT 30.000 -21.500 30.170 -20.230 ;
        RECT 30.440 -20.360 30.610 -20.230 ;
        RECT 31.890 -20.360 32.060 -20.230 ;
        RECT 30.380 -20.530 30.650 -20.360 ;
        RECT 31.850 -20.530 32.120 -20.360 ;
        RECT 30.440 -20.650 30.610 -20.530 ;
        RECT 31.890 -20.650 32.060 -20.530 ;
        RECT 30.450 -21.070 30.620 -21.030 ;
        RECT 31.870 -21.050 32.040 -21.010 ;
        RECT 32.330 -21.030 32.500 -20.230 ;
        RECT 32.900 -20.860 33.070 -19.860 ;
        RECT 33.340 -20.860 33.510 -19.860 ;
        RECT 33.780 -20.370 33.950 -19.860 ;
        RECT 34.300 -20.370 34.470 -19.860 ;
        RECT 33.720 -20.540 33.990 -20.370 ;
        RECT 34.260 -20.540 34.530 -20.370 ;
        RECT 33.780 -20.860 33.950 -20.540 ;
        RECT 34.300 -20.860 34.470 -20.540 ;
        RECT 34.740 -20.860 34.910 -19.860 ;
        RECT 35.180 -20.860 35.350 -19.860 ;
        RECT 30.370 -21.240 30.700 -21.070 ;
        RECT 31.790 -21.220 32.120 -21.050 ;
        RECT 32.330 -21.070 32.560 -21.030 ;
        RECT 30.450 -21.280 30.620 -21.240 ;
        RECT 31.870 -21.260 32.040 -21.220 ;
        RECT 32.330 -21.240 32.620 -21.070 ;
        RECT 33.500 -21.240 33.830 -21.070 ;
        RECT 34.420 -21.240 34.750 -21.070 ;
        RECT 32.330 -21.280 32.560 -21.240 ;
        RECT 27.830 -21.670 30.170 -21.500 ;
        RECT 30.000 -22.340 30.170 -21.670 ;
        RECT 30.440 -21.780 30.610 -21.500 ;
        RECT 30.420 -21.840 30.610 -21.780 ;
        RECT 31.890 -21.840 32.060 -21.500 ;
        RECT 30.380 -22.010 31.410 -21.840 ;
        RECT 31.850 -22.010 32.120 -21.840 ;
        RECT 30.420 -22.070 30.610 -22.010 ;
        RECT 30.440 -22.340 30.610 -22.070 ;
        RECT 31.890 -22.340 32.060 -22.010 ;
        RECT 32.330 -22.340 32.500 -21.280 ;
        RECT 33.580 -21.500 33.750 -21.240 ;
        RECT 35.750 -21.500 35.920 -20.230 ;
        RECT 36.190 -20.360 36.360 -20.230 ;
        RECT 37.640 -20.360 37.810 -20.230 ;
        RECT 36.130 -20.530 36.400 -20.360 ;
        RECT 37.600 -20.530 37.870 -20.360 ;
        RECT 36.190 -20.650 36.360 -20.530 ;
        RECT 37.640 -20.650 37.810 -20.530 ;
        RECT 36.200 -21.070 36.370 -21.030 ;
        RECT 37.620 -21.050 37.790 -21.010 ;
        RECT 38.080 -21.030 38.250 -20.230 ;
        RECT 38.650 -20.860 38.820 -19.860 ;
        RECT 39.090 -20.860 39.260 -19.860 ;
        RECT 39.530 -20.370 39.700 -19.860 ;
        RECT 40.050 -20.370 40.220 -19.860 ;
        RECT 39.470 -20.540 39.740 -20.370 ;
        RECT 40.010 -20.540 40.280 -20.370 ;
        RECT 39.530 -20.860 39.700 -20.540 ;
        RECT 40.050 -20.860 40.220 -20.540 ;
        RECT 40.490 -20.860 40.660 -19.860 ;
        RECT 40.930 -20.860 41.100 -19.860 ;
        RECT 36.120 -21.240 36.450 -21.070 ;
        RECT 37.540 -21.220 37.870 -21.050 ;
        RECT 38.080 -21.070 38.310 -21.030 ;
        RECT 36.200 -21.280 36.370 -21.240 ;
        RECT 37.620 -21.260 37.790 -21.220 ;
        RECT 38.080 -21.240 38.370 -21.070 ;
        RECT 39.250 -21.240 39.580 -21.070 ;
        RECT 40.170 -21.240 40.500 -21.070 ;
        RECT 38.080 -21.280 38.310 -21.240 ;
        RECT 33.580 -21.670 35.920 -21.500 ;
        RECT 35.750 -22.340 35.920 -21.670 ;
        RECT 36.190 -21.780 36.360 -21.500 ;
        RECT 36.170 -21.840 36.360 -21.780 ;
        RECT 37.640 -21.840 37.810 -21.500 ;
        RECT 36.130 -22.010 37.160 -21.840 ;
        RECT 37.600 -22.010 37.870 -21.840 ;
        RECT 36.170 -22.070 36.360 -22.010 ;
        RECT 36.190 -22.340 36.360 -22.070 ;
        RECT 37.640 -22.340 37.810 -22.010 ;
        RECT 38.080 -22.340 38.250 -21.280 ;
        RECT 39.330 -21.500 39.500 -21.240 ;
        RECT 41.500 -21.500 41.670 -20.230 ;
        RECT 41.940 -20.360 42.110 -20.230 ;
        RECT 43.390 -20.360 43.560 -20.230 ;
        RECT 41.880 -20.530 42.150 -20.360 ;
        RECT 43.350 -20.530 43.620 -20.360 ;
        RECT 41.940 -20.650 42.110 -20.530 ;
        RECT 43.390 -20.650 43.560 -20.530 ;
        RECT 41.950 -21.070 42.120 -21.030 ;
        RECT 43.370 -21.050 43.540 -21.010 ;
        RECT 43.830 -21.030 44.000 -20.230 ;
        RECT 44.400 -20.860 44.570 -19.860 ;
        RECT 44.840 -20.860 45.010 -19.860 ;
        RECT 45.280 -20.370 45.450 -19.860 ;
        RECT 45.800 -20.370 45.970 -19.860 ;
        RECT 45.220 -20.540 45.490 -20.370 ;
        RECT 45.760 -20.540 46.030 -20.370 ;
        RECT 45.280 -20.860 45.450 -20.540 ;
        RECT 45.800 -20.860 45.970 -20.540 ;
        RECT 46.240 -20.860 46.410 -19.860 ;
        RECT 46.680 -20.860 46.850 -19.860 ;
        RECT 41.870 -21.240 42.200 -21.070 ;
        RECT 43.290 -21.220 43.620 -21.050 ;
        RECT 43.830 -21.070 44.060 -21.030 ;
        RECT 41.950 -21.280 42.120 -21.240 ;
        RECT 43.370 -21.260 43.540 -21.220 ;
        RECT 43.830 -21.240 44.120 -21.070 ;
        RECT 45.000 -21.240 45.330 -21.070 ;
        RECT 45.920 -21.240 46.250 -21.070 ;
        RECT 43.830 -21.280 44.060 -21.240 ;
        RECT 39.330 -21.670 41.670 -21.500 ;
        RECT 41.500 -22.340 41.670 -21.670 ;
        RECT 41.940 -21.780 42.110 -21.500 ;
        RECT 41.920 -21.840 42.110 -21.780 ;
        RECT 43.390 -21.840 43.560 -21.500 ;
        RECT 41.880 -22.010 42.910 -21.840 ;
        RECT 43.350 -22.010 43.620 -21.840 ;
        RECT 41.920 -22.070 42.110 -22.010 ;
        RECT 41.940 -22.340 42.110 -22.070 ;
        RECT 43.390 -22.340 43.560 -22.010 ;
        RECT 43.830 -22.340 44.000 -21.280 ;
        RECT 45.080 -21.500 45.250 -21.240 ;
        RECT 47.250 -21.500 47.420 -20.230 ;
        RECT 47.690 -20.360 47.860 -20.230 ;
        RECT 49.140 -20.360 49.310 -20.230 ;
        RECT 47.630 -20.530 47.900 -20.360 ;
        RECT 49.100 -20.530 49.370 -20.360 ;
        RECT 47.690 -20.650 47.860 -20.530 ;
        RECT 49.140 -20.650 49.310 -20.530 ;
        RECT 47.700 -21.070 47.870 -21.030 ;
        RECT 49.120 -21.050 49.290 -21.010 ;
        RECT 49.580 -21.030 49.750 -20.230 ;
        RECT 50.150 -20.860 50.320 -19.860 ;
        RECT 50.590 -20.860 50.760 -19.860 ;
        RECT 51.030 -20.370 51.200 -19.860 ;
        RECT 51.550 -20.370 51.720 -19.860 ;
        RECT 50.970 -20.540 51.240 -20.370 ;
        RECT 51.510 -20.540 51.780 -20.370 ;
        RECT 51.030 -20.860 51.200 -20.540 ;
        RECT 51.550 -20.860 51.720 -20.540 ;
        RECT 51.990 -20.860 52.160 -19.860 ;
        RECT 52.430 -20.860 52.600 -19.860 ;
        RECT 47.620 -21.240 47.950 -21.070 ;
        RECT 49.040 -21.220 49.370 -21.050 ;
        RECT 49.580 -21.070 49.810 -21.030 ;
        RECT 47.700 -21.280 47.870 -21.240 ;
        RECT 49.120 -21.260 49.290 -21.220 ;
        RECT 49.580 -21.240 49.870 -21.070 ;
        RECT 50.750 -21.240 51.080 -21.070 ;
        RECT 51.670 -21.240 52.000 -21.070 ;
        RECT 49.580 -21.280 49.810 -21.240 ;
        RECT 45.080 -21.670 47.420 -21.500 ;
        RECT 47.250 -22.340 47.420 -21.670 ;
        RECT 47.690 -21.780 47.860 -21.500 ;
        RECT 47.670 -21.840 47.860 -21.780 ;
        RECT 49.140 -21.840 49.310 -21.500 ;
        RECT 47.630 -22.010 48.660 -21.840 ;
        RECT 49.100 -22.010 49.370 -21.840 ;
        RECT 47.670 -22.070 47.860 -22.010 ;
        RECT 47.690 -22.340 47.860 -22.070 ;
        RECT 49.140 -22.340 49.310 -22.010 ;
        RECT 49.580 -22.340 49.750 -21.280 ;
        RECT 50.830 -21.500 51.000 -21.240 ;
        RECT 53.000 -21.500 53.170 -20.230 ;
        RECT 53.440 -20.360 53.610 -20.230 ;
        RECT 54.890 -20.360 55.060 -20.230 ;
        RECT 53.380 -20.530 53.650 -20.360 ;
        RECT 54.850 -20.530 55.120 -20.360 ;
        RECT 53.440 -20.650 53.610 -20.530 ;
        RECT 54.890 -20.650 55.060 -20.530 ;
        RECT 53.450 -21.070 53.620 -21.030 ;
        RECT 54.870 -21.050 55.040 -21.010 ;
        RECT 55.330 -21.030 55.500 -20.230 ;
        RECT 55.900 -20.860 56.070 -19.860 ;
        RECT 56.340 -20.860 56.510 -19.860 ;
        RECT 56.780 -20.370 56.950 -19.860 ;
        RECT 57.300 -20.370 57.470 -19.860 ;
        RECT 56.720 -20.540 56.990 -20.370 ;
        RECT 57.260 -20.540 57.530 -20.370 ;
        RECT 56.780 -20.860 56.950 -20.540 ;
        RECT 57.300 -20.860 57.470 -20.540 ;
        RECT 57.740 -20.860 57.910 -19.860 ;
        RECT 58.180 -20.860 58.350 -19.860 ;
        RECT 53.370 -21.240 53.700 -21.070 ;
        RECT 54.790 -21.220 55.120 -21.050 ;
        RECT 55.330 -21.070 55.560 -21.030 ;
        RECT 53.450 -21.280 53.620 -21.240 ;
        RECT 54.870 -21.260 55.040 -21.220 ;
        RECT 55.330 -21.240 55.620 -21.070 ;
        RECT 56.500 -21.240 56.830 -21.070 ;
        RECT 57.420 -21.240 57.750 -21.070 ;
        RECT 55.330 -21.280 55.560 -21.240 ;
        RECT 50.830 -21.670 53.170 -21.500 ;
        RECT 53.000 -22.340 53.170 -21.670 ;
        RECT 53.440 -21.780 53.610 -21.500 ;
        RECT 53.420 -21.840 53.610 -21.780 ;
        RECT 54.890 -21.840 55.060 -21.500 ;
        RECT 53.380 -22.010 54.410 -21.840 ;
        RECT 54.850 -22.010 55.120 -21.840 ;
        RECT 53.420 -22.070 53.610 -22.010 ;
        RECT 53.440 -22.340 53.610 -22.070 ;
        RECT 54.890 -22.340 55.060 -22.010 ;
        RECT 55.330 -22.340 55.500 -21.280 ;
        RECT 56.580 -21.500 56.750 -21.240 ;
        RECT 58.750 -21.500 58.920 -20.230 ;
        RECT 59.190 -20.360 59.360 -20.230 ;
        RECT 60.640 -20.360 60.810 -20.230 ;
        RECT 59.130 -20.530 59.400 -20.360 ;
        RECT 60.600 -20.530 60.870 -20.360 ;
        RECT 59.190 -20.650 59.360 -20.530 ;
        RECT 60.640 -20.650 60.810 -20.530 ;
        RECT 59.200 -21.070 59.370 -21.030 ;
        RECT 60.620 -21.050 60.790 -21.010 ;
        RECT 61.080 -21.030 61.250 -20.230 ;
        RECT 61.650 -20.860 61.820 -19.860 ;
        RECT 62.090 -20.860 62.260 -19.860 ;
        RECT 62.530 -20.370 62.700 -19.860 ;
        RECT 63.050 -20.370 63.220 -19.860 ;
        RECT 62.470 -20.540 62.740 -20.370 ;
        RECT 63.010 -20.540 63.280 -20.370 ;
        RECT 62.530 -20.860 62.700 -20.540 ;
        RECT 63.050 -20.860 63.220 -20.540 ;
        RECT 63.490 -20.860 63.660 -19.860 ;
        RECT 63.930 -20.860 64.100 -19.860 ;
        RECT 59.120 -21.240 59.450 -21.070 ;
        RECT 60.540 -21.220 60.870 -21.050 ;
        RECT 61.080 -21.070 61.310 -21.030 ;
        RECT 59.200 -21.280 59.370 -21.240 ;
        RECT 60.620 -21.260 60.790 -21.220 ;
        RECT 61.080 -21.240 61.370 -21.070 ;
        RECT 62.250 -21.240 62.580 -21.070 ;
        RECT 63.170 -21.240 63.500 -21.070 ;
        RECT 61.080 -21.280 61.310 -21.240 ;
        RECT 56.580 -21.670 58.920 -21.500 ;
        RECT 58.750 -22.340 58.920 -21.670 ;
        RECT 59.190 -21.780 59.360 -21.500 ;
        RECT 59.170 -21.840 59.360 -21.780 ;
        RECT 60.640 -21.840 60.810 -21.500 ;
        RECT 59.130 -22.010 60.160 -21.840 ;
        RECT 60.600 -22.010 60.870 -21.840 ;
        RECT 59.170 -22.070 59.360 -22.010 ;
        RECT 59.190 -22.340 59.360 -22.070 ;
        RECT 60.640 -22.340 60.810 -22.010 ;
        RECT 61.080 -22.340 61.250 -21.280 ;
        RECT 62.330 -21.500 62.500 -21.240 ;
        RECT 64.500 -21.500 64.670 -20.230 ;
        RECT 64.940 -20.360 65.110 -20.230 ;
        RECT 66.390 -20.360 66.560 -20.230 ;
        RECT 64.880 -20.530 65.150 -20.360 ;
        RECT 66.350 -20.530 66.620 -20.360 ;
        RECT 64.940 -20.650 65.110 -20.530 ;
        RECT 66.390 -20.650 66.560 -20.530 ;
        RECT 64.950 -21.070 65.120 -21.030 ;
        RECT 66.370 -21.050 66.540 -21.010 ;
        RECT 66.830 -21.030 67.000 -20.230 ;
        RECT 67.400 -20.860 67.570 -19.860 ;
        RECT 67.840 -20.860 68.010 -19.860 ;
        RECT 68.280 -20.370 68.450 -19.860 ;
        RECT 68.800 -20.370 68.970 -19.860 ;
        RECT 68.220 -20.540 68.490 -20.370 ;
        RECT 68.760 -20.540 69.030 -20.370 ;
        RECT 68.280 -20.860 68.450 -20.540 ;
        RECT 68.800 -20.860 68.970 -20.540 ;
        RECT 69.240 -20.860 69.410 -19.860 ;
        RECT 69.680 -20.860 69.850 -19.860 ;
        RECT 64.870 -21.240 65.200 -21.070 ;
        RECT 66.290 -21.220 66.620 -21.050 ;
        RECT 66.830 -21.070 67.060 -21.030 ;
        RECT 64.950 -21.280 65.120 -21.240 ;
        RECT 66.370 -21.260 66.540 -21.220 ;
        RECT 66.830 -21.240 67.120 -21.070 ;
        RECT 68.000 -21.240 68.330 -21.070 ;
        RECT 68.920 -21.240 69.250 -21.070 ;
        RECT 66.830 -21.280 67.060 -21.240 ;
        RECT 62.330 -21.670 64.670 -21.500 ;
        RECT 64.500 -22.340 64.670 -21.670 ;
        RECT 64.940 -21.780 65.110 -21.500 ;
        RECT 64.920 -21.840 65.110 -21.780 ;
        RECT 66.390 -21.840 66.560 -21.500 ;
        RECT 64.880 -22.010 65.910 -21.840 ;
        RECT 66.350 -22.010 66.620 -21.840 ;
        RECT 64.920 -22.070 65.110 -22.010 ;
        RECT 64.940 -22.340 65.110 -22.070 ;
        RECT 66.390 -22.340 66.560 -22.010 ;
        RECT 66.830 -22.340 67.000 -21.280 ;
        RECT 68.080 -21.500 68.250 -21.240 ;
        RECT 70.250 -21.500 70.420 -20.230 ;
        RECT 70.690 -20.360 70.860 -20.230 ;
        RECT 72.140 -20.360 72.310 -20.230 ;
        RECT 70.630 -20.530 70.900 -20.360 ;
        RECT 72.100 -20.530 72.370 -20.360 ;
        RECT 70.690 -20.650 70.860 -20.530 ;
        RECT 72.140 -20.650 72.310 -20.530 ;
        RECT 70.700 -21.070 70.870 -21.030 ;
        RECT 72.120 -21.050 72.290 -21.010 ;
        RECT 72.580 -21.030 72.750 -20.230 ;
        RECT 73.150 -20.860 73.320 -19.860 ;
        RECT 73.590 -20.860 73.760 -19.860 ;
        RECT 74.030 -20.370 74.200 -19.860 ;
        RECT 74.550 -20.370 74.720 -19.860 ;
        RECT 73.970 -20.540 74.240 -20.370 ;
        RECT 74.510 -20.540 74.780 -20.370 ;
        RECT 74.030 -20.860 74.200 -20.540 ;
        RECT 74.550 -20.860 74.720 -20.540 ;
        RECT 74.990 -20.860 75.160 -19.860 ;
        RECT 75.430 -20.860 75.600 -19.860 ;
        RECT 70.620 -21.240 70.950 -21.070 ;
        RECT 72.040 -21.220 72.370 -21.050 ;
        RECT 72.580 -21.070 72.810 -21.030 ;
        RECT 70.700 -21.280 70.870 -21.240 ;
        RECT 72.120 -21.260 72.290 -21.220 ;
        RECT 72.580 -21.240 72.870 -21.070 ;
        RECT 73.750 -21.240 74.080 -21.070 ;
        RECT 74.670 -21.240 75.000 -21.070 ;
        RECT 72.580 -21.280 72.810 -21.240 ;
        RECT 68.080 -21.670 70.420 -21.500 ;
        RECT 70.250 -22.340 70.420 -21.670 ;
        RECT 70.690 -21.780 70.860 -21.500 ;
        RECT 70.670 -21.840 70.860 -21.780 ;
        RECT 72.140 -21.840 72.310 -21.500 ;
        RECT 70.630 -22.010 71.660 -21.840 ;
        RECT 72.100 -22.010 72.370 -21.840 ;
        RECT 70.670 -22.070 70.860 -22.010 ;
        RECT 70.690 -22.340 70.860 -22.070 ;
        RECT 72.140 -22.340 72.310 -22.010 ;
        RECT 72.580 -22.340 72.750 -21.280 ;
        RECT 73.830 -21.500 74.000 -21.240 ;
        RECT 76.000 -21.500 76.170 -20.230 ;
        RECT 76.440 -20.360 76.610 -20.230 ;
        RECT 77.890 -20.360 78.060 -20.230 ;
        RECT 76.380 -20.530 76.650 -20.360 ;
        RECT 77.850 -20.530 78.120 -20.360 ;
        RECT 76.440 -20.650 76.610 -20.530 ;
        RECT 77.890 -20.650 78.060 -20.530 ;
        RECT 76.450 -21.070 76.620 -21.030 ;
        RECT 77.870 -21.050 78.040 -21.010 ;
        RECT 78.330 -21.030 78.500 -20.230 ;
        RECT 78.900 -20.860 79.070 -19.860 ;
        RECT 79.340 -20.860 79.510 -19.860 ;
        RECT 79.780 -20.370 79.950 -19.860 ;
        RECT 80.300 -20.370 80.470 -19.860 ;
        RECT 79.720 -20.540 79.990 -20.370 ;
        RECT 80.260 -20.540 80.530 -20.370 ;
        RECT 79.780 -20.860 79.950 -20.540 ;
        RECT 80.300 -20.860 80.470 -20.540 ;
        RECT 80.740 -20.860 80.910 -19.860 ;
        RECT 81.180 -20.860 81.350 -19.860 ;
        RECT 76.370 -21.240 76.700 -21.070 ;
        RECT 77.790 -21.220 78.120 -21.050 ;
        RECT 78.330 -21.070 78.560 -21.030 ;
        RECT 76.450 -21.280 76.620 -21.240 ;
        RECT 77.870 -21.260 78.040 -21.220 ;
        RECT 78.330 -21.240 78.620 -21.070 ;
        RECT 79.500 -21.240 79.830 -21.070 ;
        RECT 80.420 -21.240 80.750 -21.070 ;
        RECT 78.330 -21.280 78.560 -21.240 ;
        RECT 73.830 -21.670 76.170 -21.500 ;
        RECT 76.000 -22.340 76.170 -21.670 ;
        RECT 76.440 -21.780 76.610 -21.500 ;
        RECT 76.420 -21.840 76.610 -21.780 ;
        RECT 77.890 -21.840 78.060 -21.500 ;
        RECT 76.380 -22.010 77.410 -21.840 ;
        RECT 77.850 -22.010 78.120 -21.840 ;
        RECT 76.420 -22.070 76.610 -22.010 ;
        RECT 76.440 -22.340 76.610 -22.070 ;
        RECT 77.890 -22.340 78.060 -22.010 ;
        RECT 78.330 -22.340 78.500 -21.280 ;
        RECT 79.580 -21.500 79.750 -21.240 ;
        RECT 81.750 -21.500 81.920 -20.230 ;
        RECT 82.190 -20.360 82.360 -20.230 ;
        RECT 83.640 -20.360 83.810 -20.230 ;
        RECT 82.130 -20.530 82.400 -20.360 ;
        RECT 83.600 -20.530 83.870 -20.360 ;
        RECT 82.190 -20.650 82.360 -20.530 ;
        RECT 83.640 -20.650 83.810 -20.530 ;
        RECT 82.200 -21.070 82.370 -21.030 ;
        RECT 83.620 -21.050 83.790 -21.010 ;
        RECT 84.080 -21.030 84.250 -20.230 ;
        RECT 84.650 -20.860 84.820 -19.860 ;
        RECT 85.090 -20.860 85.260 -19.860 ;
        RECT 85.530 -20.370 85.700 -19.860 ;
        RECT 86.050 -20.370 86.220 -19.860 ;
        RECT 85.470 -20.540 85.740 -20.370 ;
        RECT 86.010 -20.540 86.280 -20.370 ;
        RECT 85.530 -20.860 85.700 -20.540 ;
        RECT 86.050 -20.860 86.220 -20.540 ;
        RECT 86.490 -20.860 86.660 -19.860 ;
        RECT 86.930 -20.860 87.100 -19.860 ;
        RECT 82.120 -21.240 82.450 -21.070 ;
        RECT 83.540 -21.220 83.870 -21.050 ;
        RECT 84.080 -21.070 84.310 -21.030 ;
        RECT 82.200 -21.280 82.370 -21.240 ;
        RECT 83.620 -21.260 83.790 -21.220 ;
        RECT 84.080 -21.240 84.370 -21.070 ;
        RECT 85.250 -21.240 85.580 -21.070 ;
        RECT 86.170 -21.240 86.500 -21.070 ;
        RECT 84.080 -21.280 84.310 -21.240 ;
        RECT 79.580 -21.670 81.920 -21.500 ;
        RECT 81.750 -22.340 81.920 -21.670 ;
        RECT 82.190 -21.780 82.360 -21.500 ;
        RECT 82.170 -21.840 82.360 -21.780 ;
        RECT 83.640 -21.840 83.810 -21.500 ;
        RECT 82.130 -22.010 83.160 -21.840 ;
        RECT 83.600 -22.010 83.870 -21.840 ;
        RECT 82.170 -22.070 82.360 -22.010 ;
        RECT 82.190 -22.340 82.360 -22.070 ;
        RECT 83.640 -22.340 83.810 -22.010 ;
        RECT 84.080 -22.340 84.250 -21.280 ;
        RECT 85.330 -21.500 85.500 -21.240 ;
        RECT 87.500 -21.500 87.670 -20.230 ;
        RECT 87.940 -20.360 88.110 -20.230 ;
        RECT 89.390 -20.360 89.560 -20.230 ;
        RECT 87.880 -20.530 88.150 -20.360 ;
        RECT 89.350 -20.530 89.620 -20.360 ;
        RECT 87.940 -20.650 88.110 -20.530 ;
        RECT 89.390 -20.650 89.560 -20.530 ;
        RECT 87.950 -21.070 88.120 -21.030 ;
        RECT 89.370 -21.050 89.540 -21.010 ;
        RECT 89.830 -21.030 90.000 -20.230 ;
        RECT 90.400 -20.860 90.570 -19.860 ;
        RECT 90.840 -20.860 91.010 -19.860 ;
        RECT 91.280 -20.370 91.450 -19.860 ;
        RECT 91.800 -20.370 91.970 -19.860 ;
        RECT 91.220 -20.540 91.490 -20.370 ;
        RECT 91.760 -20.540 92.030 -20.370 ;
        RECT 91.280 -20.860 91.450 -20.540 ;
        RECT 91.800 -20.860 91.970 -20.540 ;
        RECT 92.240 -20.860 92.410 -19.860 ;
        RECT 92.680 -20.860 92.850 -19.860 ;
        RECT 87.870 -21.240 88.200 -21.070 ;
        RECT 89.290 -21.220 89.620 -21.050 ;
        RECT 89.830 -21.070 90.060 -21.030 ;
        RECT 87.950 -21.280 88.120 -21.240 ;
        RECT 89.370 -21.260 89.540 -21.220 ;
        RECT 89.830 -21.240 90.120 -21.070 ;
        RECT 91.000 -21.240 91.330 -21.070 ;
        RECT 91.920 -21.240 92.250 -21.070 ;
        RECT 89.830 -21.280 90.060 -21.240 ;
        RECT 85.330 -21.670 87.670 -21.500 ;
        RECT 87.500 -22.340 87.670 -21.670 ;
        RECT 87.940 -21.780 88.110 -21.500 ;
        RECT 87.920 -21.840 88.110 -21.780 ;
        RECT 89.390 -21.830 89.560 -21.500 ;
        RECT 89.040 -21.840 89.560 -21.830 ;
        RECT 87.880 -22.010 89.620 -21.840 ;
        RECT 87.920 -22.070 88.110 -22.010 ;
        RECT 87.940 -22.340 88.110 -22.070 ;
        RECT 89.390 -22.340 89.560 -22.010 ;
        RECT 89.830 -22.340 90.000 -21.280 ;
        RECT 91.080 -21.500 91.250 -21.240 ;
        RECT 93.250 -21.500 93.420 -20.230 ;
        RECT 93.690 -20.360 93.860 -20.230 ;
        RECT 93.630 -20.530 93.900 -20.360 ;
        RECT 93.690 -20.650 93.860 -20.530 ;
        RECT 93.700 -21.070 93.870 -21.030 ;
        RECT 93.620 -21.240 93.950 -21.070 ;
        RECT 93.700 -21.280 93.870 -21.240 ;
        RECT 91.080 -21.670 93.420 -21.500 ;
        RECT 93.250 -22.340 93.420 -21.670 ;
        RECT 93.690 -21.780 93.860 -21.500 ;
        RECT 93.670 -21.840 93.860 -21.780 ;
        RECT 93.630 -22.010 93.900 -21.840 ;
        RECT 93.670 -22.070 93.860 -22.010 ;
        RECT 93.690 -22.340 93.860 -22.070 ;
        RECT 5.290 -23.470 5.490 -23.440 ;
        RECT 5.180 -23.640 5.600 -23.470 ;
        RECT 6.680 -23.480 6.850 -22.800 ;
        RECT 8.170 -23.260 8.340 -23.150 ;
        RECT 8.050 -23.430 8.460 -23.260 ;
        RECT 8.170 -23.440 8.340 -23.430 ;
        RECT 9.670 -23.470 9.840 -22.800 ;
        RECT 11.050 -23.450 11.220 -23.420 ;
        RECT 11.040 -23.470 11.240 -23.450 ;
        RECT 4.640 -23.970 4.970 -23.640 ;
        RECT 6.460 -23.650 7.100 -23.480 ;
        RECT 5.310 -23.950 5.480 -23.890 ;
        RECT 4.720 -25.200 4.890 -23.970 ;
        RECT 5.180 -24.120 7.100 -23.950 ;
        RECT 7.330 -23.960 7.660 -23.630 ;
        RECT 8.870 -23.960 9.200 -23.630 ;
        RECT 9.430 -23.640 10.070 -23.470 ;
        RECT 10.930 -23.640 11.350 -23.470 ;
        RECT 16.810 -23.500 16.980 -23.470 ;
        RECT 16.790 -23.520 16.990 -23.500 ;
        RECT 18.190 -23.520 18.360 -22.800 ;
        RECT 19.660 -23.270 19.830 -23.160 ;
        RECT 19.540 -23.440 19.950 -23.270 ;
        RECT 19.660 -23.450 19.830 -23.440 ;
        RECT 21.170 -23.520 21.340 -22.800 ;
        RECT 22.550 -23.500 22.720 -23.470 ;
        RECT 28.310 -23.500 28.480 -23.470 ;
        RECT 22.540 -23.520 22.740 -23.500 ;
        RECT 28.290 -23.520 28.490 -23.500 ;
        RECT 29.690 -23.520 29.860 -22.800 ;
        RECT 31.090 -23.280 31.260 -23.170 ;
        RECT 30.970 -23.450 31.380 -23.280 ;
        RECT 31.090 -23.460 31.260 -23.450 ;
        RECT 32.670 -23.520 32.840 -22.800 ;
        RECT 34.050 -23.500 34.220 -23.470 ;
        RECT 39.810 -23.500 39.980 -23.470 ;
        RECT 34.040 -23.520 34.240 -23.500 ;
        RECT 39.790 -23.520 39.990 -23.500 ;
        RECT 41.190 -23.520 41.360 -22.800 ;
        RECT 42.660 -23.290 42.830 -23.180 ;
        RECT 42.540 -23.460 42.950 -23.290 ;
        RECT 42.660 -23.470 42.830 -23.460 ;
        RECT 44.170 -23.520 44.340 -22.800 ;
        RECT 45.550 -23.500 45.720 -23.470 ;
        RECT 51.310 -23.500 51.480 -23.470 ;
        RECT 45.540 -23.520 45.740 -23.500 ;
        RECT 51.290 -23.520 51.490 -23.500 ;
        RECT 52.690 -23.520 52.860 -22.800 ;
        RECT 54.060 -23.270 54.230 -23.160 ;
        RECT 53.940 -23.440 54.350 -23.270 ;
        RECT 54.060 -23.450 54.230 -23.440 ;
        RECT 55.670 -23.520 55.840 -22.800 ;
        RECT 57.050 -23.500 57.220 -23.470 ;
        RECT 62.810 -23.500 62.980 -23.470 ;
        RECT 57.040 -23.520 57.240 -23.500 ;
        RECT 62.790 -23.520 62.990 -23.500 ;
        RECT 64.190 -23.520 64.360 -22.800 ;
        RECT 65.740 -23.270 65.910 -23.160 ;
        RECT 65.620 -23.440 66.030 -23.270 ;
        RECT 65.740 -23.450 65.910 -23.440 ;
        RECT 67.170 -23.520 67.340 -22.800 ;
        RECT 68.550 -23.500 68.720 -23.470 ;
        RECT 74.310 -23.500 74.480 -23.470 ;
        RECT 68.540 -23.520 68.740 -23.500 ;
        RECT 74.290 -23.520 74.490 -23.500 ;
        RECT 75.690 -23.520 75.860 -22.800 ;
        RECT 77.190 -23.270 77.360 -23.160 ;
        RECT 77.070 -23.440 77.480 -23.270 ;
        RECT 77.190 -23.450 77.360 -23.440 ;
        RECT 78.670 -23.520 78.840 -22.800 ;
        RECT 80.050 -23.500 80.220 -23.470 ;
        RECT 85.810 -23.500 85.980 -23.470 ;
        RECT 80.040 -23.520 80.240 -23.500 ;
        RECT 85.790 -23.520 85.990 -23.500 ;
        RECT 87.190 -23.520 87.360 -22.800 ;
        RECT 88.760 -23.250 88.930 -23.140 ;
        RECT 88.640 -23.420 89.050 -23.250 ;
        RECT 88.760 -23.430 88.930 -23.420 ;
        RECT 90.170 -23.520 90.340 -22.800 ;
        RECT 91.550 -23.500 91.720 -23.470 ;
        RECT 91.540 -23.520 91.740 -23.500 ;
        RECT 11.040 -23.650 11.240 -23.640 ;
        RECT 11.050 -23.700 11.220 -23.650 ;
        RECT 5.310 -24.170 5.480 -24.120 ;
        RECT 6.690 -24.790 6.860 -24.120 ;
        RECT 7.410 -24.540 7.580 -23.960 ;
        RECT 8.960 -24.540 9.130 -23.960 ;
        RECT 9.430 -24.110 11.350 -23.940 ;
        RECT 11.560 -23.950 11.890 -23.620 ;
        RECT 9.680 -25.630 9.850 -24.110 ;
        RECT 11.650 -25.130 11.820 -23.950 ;
        RECT 16.140 -24.000 16.470 -23.670 ;
        RECT 16.680 -23.690 17.100 -23.520 ;
        RECT 17.960 -23.690 18.600 -23.520 ;
        RECT 16.790 -23.700 16.990 -23.690 ;
        RECT 16.810 -23.750 16.980 -23.700 ;
        RECT 16.210 -25.120 16.380 -24.000 ;
        RECT 16.680 -24.170 18.600 -24.000 ;
        RECT 18.830 -24.010 19.160 -23.680 ;
        RECT 20.370 -24.010 20.700 -23.680 ;
        RECT 20.930 -23.690 21.570 -23.520 ;
        RECT 22.430 -23.690 22.850 -23.520 ;
        RECT 22.540 -23.700 22.740 -23.690 ;
        RECT 22.550 -23.750 22.720 -23.700 ;
        RECT 23.060 -24.000 23.390 -23.670 ;
        RECT 27.640 -24.000 27.970 -23.670 ;
        RECT 28.180 -23.690 28.600 -23.520 ;
        RECT 29.460 -23.690 30.100 -23.520 ;
        RECT 28.290 -23.700 28.490 -23.690 ;
        RECT 28.310 -23.750 28.480 -23.700 ;
        RECT 30.330 -23.760 30.660 -23.680 ;
        RECT 31.870 -23.760 32.200 -23.680 ;
        RECT 32.430 -23.690 33.070 -23.520 ;
        RECT 33.930 -23.690 34.350 -23.520 ;
        RECT 34.040 -23.700 34.240 -23.690 ;
        RECT 34.050 -23.750 34.220 -23.700 ;
        RECT 30.330 -23.930 30.830 -23.760 ;
        RECT 31.700 -23.930 32.200 -23.760 ;
        RECT 18.180 -26.260 18.350 -24.170 ;
        RECT 18.910 -24.430 19.080 -24.010 ;
        RECT 20.460 -24.430 20.630 -24.010 ;
        RECT 20.930 -24.170 22.850 -24.000 ;
        RECT 21.180 -27.010 21.350 -24.170 ;
        RECT 23.140 -25.170 23.310 -24.000 ;
        RECT 27.730 -25.180 27.900 -24.000 ;
        RECT 28.180 -24.170 30.100 -24.000 ;
        RECT 30.330 -24.010 30.660 -23.930 ;
        RECT 31.870 -24.010 32.200 -23.930 ;
        RECT 34.560 -24.000 34.890 -23.670 ;
        RECT 39.140 -24.000 39.470 -23.670 ;
        RECT 39.680 -23.690 40.100 -23.520 ;
        RECT 40.960 -23.690 41.600 -23.520 ;
        RECT 39.790 -23.700 39.990 -23.690 ;
        RECT 39.810 -23.750 39.980 -23.700 ;
        RECT 41.830 -23.760 42.160 -23.680 ;
        RECT 43.370 -23.760 43.700 -23.680 ;
        RECT 43.930 -23.690 44.570 -23.520 ;
        RECT 45.430 -23.690 45.850 -23.520 ;
        RECT 45.540 -23.700 45.740 -23.690 ;
        RECT 45.550 -23.750 45.720 -23.700 ;
        RECT 41.830 -23.930 42.330 -23.760 ;
        RECT 43.200 -23.930 43.700 -23.760 ;
        RECT 29.680 -27.720 29.850 -24.170 ;
        RECT 30.410 -24.540 30.580 -24.010 ;
        RECT 31.950 -24.540 32.120 -24.010 ;
        RECT 32.430 -24.170 34.350 -24.000 ;
        RECT 32.430 -24.180 33.070 -24.170 ;
        RECT 32.680 -28.520 32.850 -24.180 ;
        RECT 34.650 -25.160 34.820 -24.000 ;
        RECT 39.230 -25.180 39.400 -24.000 ;
        RECT 39.680 -24.170 41.600 -24.000 ;
        RECT 41.830 -24.010 42.160 -23.930 ;
        RECT 43.370 -24.010 43.700 -23.930 ;
        RECT 46.060 -24.000 46.390 -23.670 ;
        RECT 50.640 -24.000 50.970 -23.670 ;
        RECT 51.180 -23.690 51.600 -23.520 ;
        RECT 52.460 -23.690 53.100 -23.520 ;
        RECT 51.290 -23.700 51.490 -23.690 ;
        RECT 51.310 -23.750 51.480 -23.700 ;
        RECT 53.330 -23.760 53.660 -23.680 ;
        RECT 54.870 -23.760 55.200 -23.680 ;
        RECT 55.430 -23.690 56.070 -23.520 ;
        RECT 56.930 -23.690 57.350 -23.520 ;
        RECT 57.040 -23.700 57.240 -23.690 ;
        RECT 57.050 -23.750 57.220 -23.700 ;
        RECT 53.330 -23.930 53.830 -23.760 ;
        RECT 54.700 -23.930 55.200 -23.760 ;
        RECT 41.180 -29.360 41.350 -24.170 ;
        RECT 41.880 -24.540 42.050 -24.010 ;
        RECT 43.470 -24.540 43.640 -24.010 ;
        RECT 43.930 -24.170 45.850 -24.000 ;
        RECT 44.180 -30.070 44.350 -24.170 ;
        RECT 46.140 -25.200 46.310 -24.000 ;
        RECT 50.720 -25.140 50.890 -24.000 ;
        RECT 51.180 -24.170 53.100 -24.000 ;
        RECT 53.330 -24.010 53.660 -23.930 ;
        RECT 54.870 -24.010 55.200 -23.930 ;
        RECT 57.560 -24.000 57.890 -23.670 ;
        RECT 62.140 -24.000 62.470 -23.670 ;
        RECT 62.680 -23.690 63.100 -23.520 ;
        RECT 63.960 -23.690 64.600 -23.520 ;
        RECT 62.790 -23.700 62.990 -23.690 ;
        RECT 62.810 -23.750 62.980 -23.700 ;
        RECT 64.830 -23.760 65.160 -23.680 ;
        RECT 66.370 -23.760 66.700 -23.680 ;
        RECT 66.930 -23.690 67.570 -23.520 ;
        RECT 68.430 -23.690 68.850 -23.520 ;
        RECT 68.540 -23.700 68.740 -23.690 ;
        RECT 68.550 -23.750 68.720 -23.700 ;
        RECT 64.830 -23.930 65.330 -23.760 ;
        RECT 66.200 -23.930 66.700 -23.760 ;
        RECT 52.680 -30.250 52.850 -24.170 ;
        RECT 53.400 -24.540 53.570 -24.010 ;
        RECT 54.950 -24.540 55.120 -24.010 ;
        RECT 55.430 -24.170 57.350 -24.000 ;
        RECT 55.680 -29.380 55.850 -24.170 ;
        RECT 57.650 -25.160 57.820 -24.000 ;
        RECT 62.220 -25.120 62.390 -24.000 ;
        RECT 62.680 -24.170 64.600 -24.000 ;
        RECT 64.830 -24.010 65.160 -23.930 ;
        RECT 66.370 -24.010 66.700 -23.930 ;
        RECT 69.060 -24.000 69.390 -23.670 ;
        RECT 73.640 -24.000 73.970 -23.670 ;
        RECT 74.180 -23.690 74.600 -23.520 ;
        RECT 75.460 -23.690 76.100 -23.520 ;
        RECT 74.290 -23.700 74.490 -23.690 ;
        RECT 74.310 -23.750 74.480 -23.700 ;
        RECT 76.330 -23.760 76.660 -23.680 ;
        RECT 77.870 -23.760 78.200 -23.680 ;
        RECT 78.430 -23.690 79.070 -23.520 ;
        RECT 79.930 -23.690 80.350 -23.520 ;
        RECT 80.040 -23.700 80.240 -23.690 ;
        RECT 80.050 -23.750 80.220 -23.700 ;
        RECT 76.330 -23.930 76.830 -23.760 ;
        RECT 77.700 -23.930 78.200 -23.760 ;
        RECT 64.180 -28.580 64.350 -24.170 ;
        RECT 64.910 -24.540 65.080 -24.010 ;
        RECT 66.440 -24.540 66.610 -24.010 ;
        RECT 66.930 -24.170 68.850 -24.000 ;
        RECT 67.180 -27.860 67.350 -24.170 ;
        RECT 69.140 -25.160 69.310 -24.000 ;
        RECT 73.720 -25.160 73.890 -24.000 ;
        RECT 74.180 -24.170 76.100 -24.000 ;
        RECT 76.330 -24.010 76.660 -23.930 ;
        RECT 77.870 -24.010 78.200 -23.930 ;
        RECT 80.560 -24.000 80.890 -23.670 ;
        RECT 85.140 -24.000 85.470 -23.670 ;
        RECT 85.680 -23.690 86.100 -23.520 ;
        RECT 86.960 -23.690 87.600 -23.520 ;
        RECT 85.790 -23.700 85.990 -23.690 ;
        RECT 85.810 -23.750 85.980 -23.700 ;
        RECT 87.830 -23.760 88.160 -23.680 ;
        RECT 89.370 -23.760 89.700 -23.680 ;
        RECT 89.930 -23.690 90.570 -23.520 ;
        RECT 91.430 -23.690 91.850 -23.520 ;
        RECT 91.540 -23.700 91.740 -23.690 ;
        RECT 91.550 -23.750 91.720 -23.700 ;
        RECT 87.830 -23.930 88.330 -23.760 ;
        RECT 89.200 -23.930 89.700 -23.760 ;
        RECT 75.680 -27.230 75.850 -24.170 ;
        RECT 76.420 -24.540 76.590 -24.010 ;
        RECT 77.950 -24.540 78.120 -24.010 ;
        RECT 78.430 -24.170 80.350 -24.000 ;
        RECT 78.680 -26.600 78.850 -24.170 ;
        RECT 80.640 -25.190 80.810 -24.000 ;
        RECT 85.220 -25.170 85.390 -24.000 ;
        RECT 85.680 -24.170 87.600 -24.000 ;
        RECT 87.830 -24.010 88.160 -23.930 ;
        RECT 89.370 -24.010 89.700 -23.930 ;
        RECT 92.060 -24.000 92.390 -23.670 ;
        RECT 87.180 -26.100 87.350 -24.170 ;
        RECT 87.910 -24.540 88.080 -24.010 ;
        RECT 89.430 -24.540 89.600 -24.010 ;
        RECT 89.930 -24.170 91.850 -24.000 ;
        RECT 90.180 -25.600 90.350 -24.170 ;
        RECT 92.160 -24.870 92.330 -24.000 ;
        RECT 92.060 -25.210 92.360 -24.870 ;
        RECT -37.290 -31.460 -36.960 -31.290 ;
        RECT -33.240 -31.460 -32.910 -31.290 ;
        RECT -25.790 -31.460 -25.460 -31.290 ;
        RECT -21.740 -31.460 -21.410 -31.290 ;
        RECT -13.970 -31.460 -13.640 -31.290 ;
        RECT -9.920 -31.460 -9.590 -31.290 ;
        RECT -2.160 -31.460 -1.830 -31.290 ;
        RECT 1.890 -31.460 2.220 -31.290 ;
        RECT 9.650 -31.460 9.980 -31.290 ;
        RECT 13.700 -31.460 14.030 -31.290 ;
        RECT 21.470 -31.460 21.800 -31.290 ;
        RECT 25.520 -31.460 25.850 -31.290 ;
        RECT 33.290 -31.460 33.620 -31.290 ;
        RECT 37.340 -31.460 37.670 -31.290 ;
        RECT 45.110 -31.460 45.440 -31.290 ;
        RECT 49.160 -31.460 49.490 -31.290 ;
        RECT 56.930 -31.460 57.260 -31.290 ;
        RECT 60.980 -31.460 61.310 -31.290 ;
        RECT 68.750 -31.460 69.080 -31.290 ;
        RECT 72.800 -31.460 73.130 -31.290 ;
        RECT 80.570 -31.460 80.900 -31.290 ;
        RECT 84.620 -31.460 84.950 -31.290 ;
        RECT 92.410 -31.460 92.740 -31.290 ;
        RECT 96.460 -31.460 96.790 -31.290 ;
        RECT 104.250 -31.460 104.580 -31.290 ;
        RECT 108.300 -31.460 108.630 -31.290 ;
        RECT 116.120 -31.460 116.450 -31.290 ;
        RECT 120.170 -31.460 120.500 -31.290 ;
        RECT 127.990 -31.460 128.320 -31.290 ;
        RECT 132.040 -31.460 132.370 -31.290 ;
        RECT 137.000 -31.460 137.330 -31.290 ;
        RECT 141.050 -31.460 141.380 -31.290 ;
        RECT -37.440 -35.890 -37.270 -31.710 ;
        RECT -37.000 -33.660 -36.830 -31.710 ;
        RECT -37.000 -33.830 -36.790 -33.660 ;
        RECT -37.000 -35.280 -36.830 -33.830 ;
        RECT -37.000 -35.450 -36.790 -35.280 ;
        RECT -37.000 -35.710 -36.830 -35.450 ;
        RECT -35.880 -35.890 -35.710 -31.710 ;
        RECT -35.440 -33.650 -35.270 -31.710 ;
        RECT -34.910 -33.650 -34.740 -31.710 ;
        RECT -35.440 -33.820 -34.740 -33.650 ;
        RECT -35.440 -35.270 -35.270 -33.820 ;
        RECT -34.910 -35.270 -34.740 -33.820 ;
        RECT -35.440 -35.440 -35.250 -35.270 ;
        RECT -34.930 -35.440 -34.740 -35.270 ;
        RECT -35.440 -35.710 -35.270 -35.440 ;
        RECT -34.910 -35.710 -34.740 -35.440 ;
        RECT -37.440 -36.060 -35.710 -35.890 ;
        RECT -34.470 -35.890 -34.300 -31.710 ;
        RECT -33.380 -33.630 -33.210 -31.710 ;
        RECT -33.420 -33.800 -33.210 -33.630 ;
        RECT -33.380 -35.280 -33.210 -33.800 ;
        RECT -33.420 -35.450 -33.210 -35.280 ;
        RECT -33.380 -35.710 -33.210 -35.450 ;
        RECT -32.940 -35.890 -32.770 -31.710 ;
        RECT -32.290 -33.930 -32.120 -33.520 ;
        RECT -34.470 -35.950 -32.770 -35.890 ;
        RECT -35.880 -36.290 -35.710 -36.060 ;
        RECT -35.530 -36.060 -32.770 -35.950 ;
        RECT -25.940 -35.890 -25.770 -31.710 ;
        RECT -25.500 -33.660 -25.330 -31.710 ;
        RECT -25.500 -33.830 -25.290 -33.660 ;
        RECT -25.500 -35.280 -25.330 -33.830 ;
        RECT -25.500 -35.450 -25.290 -35.280 ;
        RECT -25.500 -35.710 -25.330 -35.450 ;
        RECT -24.380 -35.890 -24.210 -31.710 ;
        RECT -23.940 -33.650 -23.770 -31.710 ;
        RECT -23.410 -33.650 -23.240 -31.710 ;
        RECT -23.940 -33.820 -23.240 -33.650 ;
        RECT -23.940 -35.270 -23.770 -33.820 ;
        RECT -23.410 -35.270 -23.240 -33.820 ;
        RECT -23.940 -35.440 -23.750 -35.270 ;
        RECT -23.430 -35.440 -23.240 -35.270 ;
        RECT -23.940 -35.710 -23.770 -35.440 ;
        RECT -23.410 -35.710 -23.240 -35.440 ;
        RECT -25.940 -36.060 -24.210 -35.890 ;
        RECT -22.970 -35.890 -22.800 -31.710 ;
        RECT -21.880 -33.630 -21.710 -31.710 ;
        RECT -21.920 -33.800 -21.710 -33.630 ;
        RECT -21.880 -35.280 -21.710 -33.800 ;
        RECT -21.920 -35.450 -21.710 -35.280 ;
        RECT -21.880 -35.710 -21.710 -35.450 ;
        RECT -21.440 -35.890 -21.270 -31.710 ;
        RECT -20.790 -33.930 -20.620 -33.520 ;
        RECT -22.970 -35.950 -21.270 -35.890 ;
        RECT -35.530 -36.120 -34.300 -36.060 ;
        RECT -36.790 -36.500 -36.460 -36.330 ;
        RECT -35.880 -36.460 -34.640 -36.290 ;
        RECT -37.830 -36.970 -37.660 -36.640 ;
        RECT -37.880 -37.700 -37.710 -37.150 ;
        RECT -38.230 -41.160 -38.060 -39.160 ;
        RECT -38.230 -41.550 -37.670 -41.380 ;
        RECT -38.230 -43.780 -38.060 -41.550 ;
        RECT -37.440 -43.780 -37.270 -37.150 ;
        RECT -37.830 -44.240 -37.660 -43.910 ;
        RECT -36.840 -44.700 -36.670 -36.700 ;
        RECT -36.400 -44.700 -36.230 -36.700 ;
        RECT -35.880 -44.700 -35.710 -36.460 ;
        RECT -35.440 -44.700 -35.270 -36.700 ;
        RECT -34.910 -44.700 -34.740 -36.700 ;
        RECT -34.470 -44.700 -34.300 -36.120 ;
        RECT -24.380 -36.290 -24.210 -36.060 ;
        RECT -24.030 -36.060 -21.270 -35.950 ;
        RECT -14.120 -35.890 -13.950 -31.710 ;
        RECT -13.680 -33.660 -13.510 -31.710 ;
        RECT -13.680 -33.830 -13.470 -33.660 ;
        RECT -13.680 -35.280 -13.510 -33.830 ;
        RECT -13.680 -35.450 -13.470 -35.280 ;
        RECT -13.680 -35.710 -13.510 -35.450 ;
        RECT -12.560 -35.890 -12.390 -31.710 ;
        RECT -12.120 -33.650 -11.950 -31.710 ;
        RECT -11.590 -33.650 -11.420 -31.710 ;
        RECT -12.120 -33.820 -11.420 -33.650 ;
        RECT -12.120 -35.270 -11.950 -33.820 ;
        RECT -11.590 -35.270 -11.420 -33.820 ;
        RECT -12.120 -35.440 -11.930 -35.270 ;
        RECT -11.610 -35.440 -11.420 -35.270 ;
        RECT -12.120 -35.710 -11.950 -35.440 ;
        RECT -11.590 -35.710 -11.420 -35.440 ;
        RECT -14.120 -36.060 -12.390 -35.890 ;
        RECT -11.150 -35.890 -10.980 -31.710 ;
        RECT -10.060 -33.630 -9.890 -31.710 ;
        RECT -10.100 -33.800 -9.890 -33.630 ;
        RECT -10.060 -35.280 -9.890 -33.800 ;
        RECT -10.100 -35.450 -9.890 -35.280 ;
        RECT -10.060 -35.710 -9.890 -35.450 ;
        RECT -9.620 -35.890 -9.450 -31.710 ;
        RECT -8.970 -33.930 -8.800 -33.520 ;
        RECT -11.150 -35.950 -9.450 -35.890 ;
        RECT -24.030 -36.120 -22.800 -36.060 ;
        RECT -33.720 -36.490 -33.390 -36.320 ;
        RECT -25.290 -36.500 -24.960 -36.330 ;
        RECT -24.380 -36.460 -23.140 -36.290 ;
        RECT -33.950 -44.700 -33.780 -36.700 ;
        RECT -33.510 -44.700 -33.340 -36.700 ;
        RECT -32.550 -36.980 -32.380 -36.650 ;
        RECT -26.330 -36.970 -26.160 -36.640 ;
        RECT -32.940 -41.140 -32.770 -37.150 ;
        RECT -32.500 -37.700 -32.330 -37.150 ;
        RECT -26.380 -37.700 -26.210 -37.150 ;
        RECT -32.150 -41.140 -31.980 -39.140 ;
        RECT -26.730 -41.160 -26.560 -39.160 ;
        RECT -32.500 -44.170 -32.330 -41.280 ;
        RECT -26.730 -41.550 -26.170 -41.380 ;
        RECT -26.730 -43.780 -26.560 -41.550 ;
        RECT -25.940 -43.780 -25.770 -37.150 ;
        RECT -32.500 -44.340 -31.980 -44.170 ;
        RECT -26.330 -44.240 -26.160 -43.910 ;
        RECT -32.150 -44.680 -31.980 -44.340 ;
        RECT -25.340 -44.700 -25.170 -36.700 ;
        RECT -24.900 -44.700 -24.730 -36.700 ;
        RECT -24.380 -44.700 -24.210 -36.460 ;
        RECT -23.940 -44.700 -23.770 -36.700 ;
        RECT -23.410 -44.700 -23.240 -36.700 ;
        RECT -22.970 -44.700 -22.800 -36.120 ;
        RECT -12.560 -36.290 -12.390 -36.060 ;
        RECT -12.210 -36.060 -9.450 -35.950 ;
        RECT -2.310 -35.890 -2.140 -31.710 ;
        RECT -1.870 -33.660 -1.700 -31.710 ;
        RECT -1.870 -33.830 -1.660 -33.660 ;
        RECT -1.870 -35.280 -1.700 -33.830 ;
        RECT -1.870 -35.450 -1.660 -35.280 ;
        RECT -1.870 -35.710 -1.700 -35.450 ;
        RECT -0.750 -35.890 -0.580 -31.710 ;
        RECT -0.310 -33.650 -0.140 -31.710 ;
        RECT 0.220 -33.650 0.390 -31.710 ;
        RECT -0.310 -33.820 0.390 -33.650 ;
        RECT -0.310 -35.270 -0.140 -33.820 ;
        RECT 0.220 -35.270 0.390 -33.820 ;
        RECT -0.310 -35.440 -0.120 -35.270 ;
        RECT 0.200 -35.440 0.390 -35.270 ;
        RECT -0.310 -35.710 -0.140 -35.440 ;
        RECT 0.220 -35.710 0.390 -35.440 ;
        RECT -2.310 -36.060 -0.580 -35.890 ;
        RECT 0.660 -35.890 0.830 -31.710 ;
        RECT 1.750 -33.630 1.920 -31.710 ;
        RECT 1.710 -33.800 1.920 -33.630 ;
        RECT 1.750 -35.280 1.920 -33.800 ;
        RECT 1.710 -35.450 1.920 -35.280 ;
        RECT 1.750 -35.710 1.920 -35.450 ;
        RECT 2.190 -35.890 2.360 -31.710 ;
        RECT 2.840 -33.930 3.010 -33.520 ;
        RECT 0.660 -35.950 2.360 -35.890 ;
        RECT -12.210 -36.120 -10.980 -36.060 ;
        RECT -22.220 -36.490 -21.890 -36.320 ;
        RECT -13.470 -36.500 -13.140 -36.330 ;
        RECT -12.560 -36.460 -11.320 -36.290 ;
        RECT -22.450 -44.700 -22.280 -36.700 ;
        RECT -22.010 -44.700 -21.840 -36.700 ;
        RECT -21.050 -36.980 -20.880 -36.650 ;
        RECT -14.510 -36.970 -14.340 -36.640 ;
        RECT -21.440 -41.140 -21.270 -37.150 ;
        RECT -21.000 -37.700 -20.830 -37.150 ;
        RECT -14.560 -37.700 -14.390 -37.150 ;
        RECT -20.650 -41.140 -20.480 -39.140 ;
        RECT -14.910 -41.160 -14.740 -39.160 ;
        RECT -21.000 -44.170 -20.830 -41.280 ;
        RECT -14.910 -41.550 -14.350 -41.380 ;
        RECT -14.910 -43.780 -14.740 -41.550 ;
        RECT -14.120 -43.780 -13.950 -37.150 ;
        RECT -21.000 -44.340 -20.480 -44.170 ;
        RECT -14.510 -44.240 -14.340 -43.910 ;
        RECT -20.650 -44.670 -20.480 -44.340 ;
        RECT -13.520 -44.700 -13.350 -36.700 ;
        RECT -13.080 -44.700 -12.910 -36.700 ;
        RECT -12.560 -44.700 -12.390 -36.460 ;
        RECT -12.120 -44.700 -11.950 -36.700 ;
        RECT -11.590 -44.700 -11.420 -36.700 ;
        RECT -11.150 -44.700 -10.980 -36.120 ;
        RECT -0.750 -36.290 -0.580 -36.060 ;
        RECT -0.400 -36.060 2.360 -35.950 ;
        RECT 9.500 -35.890 9.670 -31.710 ;
        RECT 9.940 -33.660 10.110 -31.710 ;
        RECT 9.940 -33.830 10.150 -33.660 ;
        RECT 9.940 -35.280 10.110 -33.830 ;
        RECT 9.940 -35.450 10.150 -35.280 ;
        RECT 9.940 -35.710 10.110 -35.450 ;
        RECT 11.060 -35.890 11.230 -31.710 ;
        RECT 11.500 -33.650 11.670 -31.710 ;
        RECT 12.030 -33.650 12.200 -31.710 ;
        RECT 11.500 -33.820 12.200 -33.650 ;
        RECT 11.500 -35.270 11.670 -33.820 ;
        RECT 12.030 -35.270 12.200 -33.820 ;
        RECT 11.500 -35.440 11.690 -35.270 ;
        RECT 12.010 -35.440 12.200 -35.270 ;
        RECT 11.500 -35.710 11.670 -35.440 ;
        RECT 12.030 -35.710 12.200 -35.440 ;
        RECT 9.500 -36.060 11.230 -35.890 ;
        RECT 12.470 -35.890 12.640 -31.710 ;
        RECT 13.560 -33.630 13.730 -31.710 ;
        RECT 13.520 -33.800 13.730 -33.630 ;
        RECT 13.560 -35.280 13.730 -33.800 ;
        RECT 13.520 -35.450 13.730 -35.280 ;
        RECT 13.560 -35.710 13.730 -35.450 ;
        RECT 14.000 -35.890 14.170 -31.710 ;
        RECT 14.650 -33.930 14.820 -33.520 ;
        RECT 12.470 -35.950 14.170 -35.890 ;
        RECT -0.400 -36.120 0.830 -36.060 ;
        RECT -10.400 -36.490 -10.070 -36.320 ;
        RECT -1.660 -36.500 -1.330 -36.330 ;
        RECT -0.750 -36.460 0.490 -36.290 ;
        RECT -10.630 -44.700 -10.460 -36.700 ;
        RECT -10.190 -44.700 -10.020 -36.700 ;
        RECT -9.230 -36.980 -9.060 -36.650 ;
        RECT -2.700 -36.970 -2.530 -36.640 ;
        RECT -9.620 -41.140 -9.450 -37.150 ;
        RECT -9.180 -37.700 -9.010 -37.150 ;
        RECT -2.750 -37.700 -2.580 -37.150 ;
        RECT -8.830 -41.140 -8.660 -39.140 ;
        RECT -3.100 -41.160 -2.930 -39.160 ;
        RECT -9.180 -44.170 -9.010 -41.280 ;
        RECT -3.100 -41.550 -2.540 -41.380 ;
        RECT -3.100 -43.780 -2.930 -41.550 ;
        RECT -2.310 -43.780 -2.140 -37.150 ;
        RECT -9.180 -44.340 -8.660 -44.170 ;
        RECT -2.700 -44.240 -2.530 -43.910 ;
        RECT -8.830 -44.670 -8.660 -44.340 ;
        RECT -1.710 -44.700 -1.540 -36.700 ;
        RECT -1.270 -44.700 -1.100 -36.700 ;
        RECT -0.750 -44.700 -0.580 -36.460 ;
        RECT -0.310 -44.700 -0.140 -36.700 ;
        RECT 0.220 -44.700 0.390 -36.700 ;
        RECT 0.660 -44.700 0.830 -36.120 ;
        RECT 11.060 -36.290 11.230 -36.060 ;
        RECT 11.410 -36.060 14.170 -35.950 ;
        RECT 21.320 -35.890 21.490 -31.710 ;
        RECT 21.760 -33.660 21.930 -31.710 ;
        RECT 21.760 -33.830 21.970 -33.660 ;
        RECT 21.760 -35.280 21.930 -33.830 ;
        RECT 21.760 -35.450 21.970 -35.280 ;
        RECT 21.760 -35.710 21.930 -35.450 ;
        RECT 22.880 -35.890 23.050 -31.710 ;
        RECT 23.320 -33.650 23.490 -31.710 ;
        RECT 23.850 -33.650 24.020 -31.710 ;
        RECT 23.320 -33.820 24.020 -33.650 ;
        RECT 23.320 -35.270 23.490 -33.820 ;
        RECT 23.850 -35.270 24.020 -33.820 ;
        RECT 23.320 -35.440 23.510 -35.270 ;
        RECT 23.830 -35.440 24.020 -35.270 ;
        RECT 23.320 -35.710 23.490 -35.440 ;
        RECT 23.850 -35.710 24.020 -35.440 ;
        RECT 21.320 -36.060 23.050 -35.890 ;
        RECT 24.290 -35.890 24.460 -31.710 ;
        RECT 25.380 -33.630 25.550 -31.710 ;
        RECT 25.340 -33.800 25.550 -33.630 ;
        RECT 25.380 -35.280 25.550 -33.800 ;
        RECT 25.340 -35.450 25.550 -35.280 ;
        RECT 25.380 -35.710 25.550 -35.450 ;
        RECT 25.820 -35.890 25.990 -31.710 ;
        RECT 26.470 -33.930 26.640 -33.520 ;
        RECT 24.290 -35.950 25.990 -35.890 ;
        RECT 11.410 -36.120 12.640 -36.060 ;
        RECT 1.410 -36.490 1.740 -36.320 ;
        RECT 10.150 -36.500 10.480 -36.330 ;
        RECT 11.060 -36.460 12.300 -36.290 ;
        RECT 1.180 -44.700 1.350 -36.700 ;
        RECT 1.620 -44.700 1.790 -36.700 ;
        RECT 2.580 -36.980 2.750 -36.650 ;
        RECT 9.110 -36.970 9.280 -36.640 ;
        RECT 2.190 -41.140 2.360 -37.150 ;
        RECT 2.630 -37.700 2.800 -37.150 ;
        RECT 9.060 -37.700 9.230 -37.150 ;
        RECT 2.980 -41.140 3.150 -39.140 ;
        RECT 8.710 -41.160 8.880 -39.160 ;
        RECT 2.630 -44.170 2.800 -41.280 ;
        RECT 8.710 -41.550 9.270 -41.380 ;
        RECT 8.710 -43.780 8.880 -41.550 ;
        RECT 9.500 -43.780 9.670 -37.150 ;
        RECT 2.630 -44.340 3.150 -44.170 ;
        RECT 9.110 -44.240 9.280 -43.910 ;
        RECT 2.980 -44.670 3.150 -44.340 ;
        RECT 10.100 -44.700 10.270 -36.700 ;
        RECT 10.540 -44.700 10.710 -36.700 ;
        RECT 11.060 -44.700 11.230 -36.460 ;
        RECT 11.500 -44.700 11.670 -36.700 ;
        RECT 12.030 -44.700 12.200 -36.700 ;
        RECT 12.470 -44.700 12.640 -36.120 ;
        RECT 22.880 -36.290 23.050 -36.060 ;
        RECT 23.230 -36.060 25.990 -35.950 ;
        RECT 33.140 -35.890 33.310 -31.710 ;
        RECT 33.580 -33.660 33.750 -31.710 ;
        RECT 33.580 -33.830 33.790 -33.660 ;
        RECT 33.580 -35.280 33.750 -33.830 ;
        RECT 33.580 -35.450 33.790 -35.280 ;
        RECT 33.580 -35.710 33.750 -35.450 ;
        RECT 34.700 -35.890 34.870 -31.710 ;
        RECT 35.140 -33.650 35.310 -31.710 ;
        RECT 35.670 -33.650 35.840 -31.710 ;
        RECT 35.140 -33.820 35.840 -33.650 ;
        RECT 35.140 -35.270 35.310 -33.820 ;
        RECT 35.670 -35.270 35.840 -33.820 ;
        RECT 35.140 -35.440 35.330 -35.270 ;
        RECT 35.650 -35.440 35.840 -35.270 ;
        RECT 35.140 -35.710 35.310 -35.440 ;
        RECT 35.670 -35.710 35.840 -35.440 ;
        RECT 33.140 -36.060 34.870 -35.890 ;
        RECT 36.110 -35.890 36.280 -31.710 ;
        RECT 37.200 -33.630 37.370 -31.710 ;
        RECT 37.160 -33.800 37.370 -33.630 ;
        RECT 37.200 -35.280 37.370 -33.800 ;
        RECT 37.160 -35.450 37.370 -35.280 ;
        RECT 37.200 -35.710 37.370 -35.450 ;
        RECT 37.640 -35.890 37.810 -31.710 ;
        RECT 38.290 -33.930 38.460 -33.520 ;
        RECT 36.110 -35.950 37.810 -35.890 ;
        RECT 23.230 -36.120 24.460 -36.060 ;
        RECT 13.220 -36.490 13.550 -36.320 ;
        RECT 21.970 -36.500 22.300 -36.330 ;
        RECT 22.880 -36.460 24.120 -36.290 ;
        RECT 12.990 -44.700 13.160 -36.700 ;
        RECT 13.430 -44.700 13.600 -36.700 ;
        RECT 14.390 -36.980 14.560 -36.650 ;
        RECT 20.930 -36.970 21.100 -36.640 ;
        RECT 14.000 -41.140 14.170 -37.150 ;
        RECT 14.440 -37.700 14.610 -37.150 ;
        RECT 20.880 -37.700 21.050 -37.150 ;
        RECT 14.790 -41.140 14.960 -39.140 ;
        RECT 20.530 -41.160 20.700 -39.160 ;
        RECT 14.440 -44.170 14.610 -41.280 ;
        RECT 20.530 -41.550 21.090 -41.380 ;
        RECT 20.530 -43.780 20.700 -41.550 ;
        RECT 21.320 -43.780 21.490 -37.150 ;
        RECT 14.440 -44.340 14.960 -44.170 ;
        RECT 20.930 -44.240 21.100 -43.910 ;
        RECT 14.790 -44.670 14.960 -44.340 ;
        RECT 21.920 -44.700 22.090 -36.700 ;
        RECT 22.360 -44.700 22.530 -36.700 ;
        RECT 22.880 -44.700 23.050 -36.460 ;
        RECT 23.320 -44.700 23.490 -36.700 ;
        RECT 23.850 -44.700 24.020 -36.700 ;
        RECT 24.290 -44.700 24.460 -36.120 ;
        RECT 34.700 -36.290 34.870 -36.060 ;
        RECT 35.050 -36.060 37.810 -35.950 ;
        RECT 44.960 -35.890 45.130 -31.710 ;
        RECT 45.400 -33.660 45.570 -31.710 ;
        RECT 45.400 -33.830 45.610 -33.660 ;
        RECT 45.400 -35.280 45.570 -33.830 ;
        RECT 45.400 -35.450 45.610 -35.280 ;
        RECT 45.400 -35.710 45.570 -35.450 ;
        RECT 46.520 -35.890 46.690 -31.710 ;
        RECT 46.960 -33.650 47.130 -31.710 ;
        RECT 47.490 -33.650 47.660 -31.710 ;
        RECT 46.960 -33.820 47.660 -33.650 ;
        RECT 46.960 -35.270 47.130 -33.820 ;
        RECT 47.490 -35.270 47.660 -33.820 ;
        RECT 46.960 -35.440 47.150 -35.270 ;
        RECT 47.470 -35.440 47.660 -35.270 ;
        RECT 46.960 -35.710 47.130 -35.440 ;
        RECT 47.490 -35.710 47.660 -35.440 ;
        RECT 44.960 -36.060 46.690 -35.890 ;
        RECT 47.930 -35.890 48.100 -31.710 ;
        RECT 49.020 -33.630 49.190 -31.710 ;
        RECT 48.980 -33.800 49.190 -33.630 ;
        RECT 49.020 -35.280 49.190 -33.800 ;
        RECT 48.980 -35.450 49.190 -35.280 ;
        RECT 49.020 -35.710 49.190 -35.450 ;
        RECT 49.460 -35.890 49.630 -31.710 ;
        RECT 50.110 -33.930 50.280 -33.520 ;
        RECT 47.930 -35.950 49.630 -35.890 ;
        RECT 35.050 -36.120 36.280 -36.060 ;
        RECT 25.040 -36.490 25.370 -36.320 ;
        RECT 33.790 -36.500 34.120 -36.330 ;
        RECT 34.700 -36.460 35.940 -36.290 ;
        RECT 24.810 -44.700 24.980 -36.700 ;
        RECT 25.250 -44.700 25.420 -36.700 ;
        RECT 26.210 -36.980 26.380 -36.650 ;
        RECT 32.750 -36.970 32.920 -36.640 ;
        RECT 25.820 -41.140 25.990 -37.150 ;
        RECT 26.260 -37.700 26.430 -37.150 ;
        RECT 32.700 -37.700 32.870 -37.150 ;
        RECT 26.610 -41.140 26.780 -39.140 ;
        RECT 32.350 -41.160 32.520 -39.160 ;
        RECT 26.260 -44.170 26.430 -41.280 ;
        RECT 32.350 -41.550 32.910 -41.380 ;
        RECT 32.350 -43.780 32.520 -41.550 ;
        RECT 33.140 -43.780 33.310 -37.150 ;
        RECT 26.260 -44.340 26.780 -44.170 ;
        RECT 32.750 -44.240 32.920 -43.910 ;
        RECT 26.610 -44.670 26.780 -44.340 ;
        RECT 33.740 -44.700 33.910 -36.700 ;
        RECT 34.180 -44.700 34.350 -36.700 ;
        RECT 34.700 -44.700 34.870 -36.460 ;
        RECT 35.140 -44.700 35.310 -36.700 ;
        RECT 35.670 -44.700 35.840 -36.700 ;
        RECT 36.110 -44.700 36.280 -36.120 ;
        RECT 46.520 -36.290 46.690 -36.060 ;
        RECT 46.870 -36.060 49.630 -35.950 ;
        RECT 56.780 -35.890 56.950 -31.710 ;
        RECT 57.220 -33.660 57.390 -31.710 ;
        RECT 57.220 -33.830 57.430 -33.660 ;
        RECT 57.220 -35.280 57.390 -33.830 ;
        RECT 57.220 -35.450 57.430 -35.280 ;
        RECT 57.220 -35.710 57.390 -35.450 ;
        RECT 58.340 -35.890 58.510 -31.710 ;
        RECT 58.780 -33.650 58.950 -31.710 ;
        RECT 59.310 -33.650 59.480 -31.710 ;
        RECT 58.780 -33.820 59.480 -33.650 ;
        RECT 58.780 -35.270 58.950 -33.820 ;
        RECT 59.310 -35.270 59.480 -33.820 ;
        RECT 58.780 -35.440 58.970 -35.270 ;
        RECT 59.290 -35.440 59.480 -35.270 ;
        RECT 58.780 -35.710 58.950 -35.440 ;
        RECT 59.310 -35.710 59.480 -35.440 ;
        RECT 56.780 -36.060 58.510 -35.890 ;
        RECT 59.750 -35.890 59.920 -31.710 ;
        RECT 60.840 -33.630 61.010 -31.710 ;
        RECT 60.800 -33.800 61.010 -33.630 ;
        RECT 60.840 -35.280 61.010 -33.800 ;
        RECT 60.800 -35.450 61.010 -35.280 ;
        RECT 60.840 -35.710 61.010 -35.450 ;
        RECT 61.280 -35.890 61.450 -31.710 ;
        RECT 61.930 -33.930 62.100 -33.520 ;
        RECT 59.750 -35.950 61.450 -35.890 ;
        RECT 46.870 -36.120 48.100 -36.060 ;
        RECT 36.860 -36.490 37.190 -36.320 ;
        RECT 45.610 -36.500 45.940 -36.330 ;
        RECT 46.520 -36.460 47.760 -36.290 ;
        RECT 36.630 -44.700 36.800 -36.700 ;
        RECT 37.070 -44.700 37.240 -36.700 ;
        RECT 38.030 -36.980 38.200 -36.650 ;
        RECT 44.570 -36.970 44.740 -36.640 ;
        RECT 37.640 -41.140 37.810 -37.150 ;
        RECT 38.080 -37.700 38.250 -37.150 ;
        RECT 44.520 -37.700 44.690 -37.150 ;
        RECT 38.430 -41.140 38.600 -39.140 ;
        RECT 44.170 -41.160 44.340 -39.160 ;
        RECT 38.080 -44.170 38.250 -41.280 ;
        RECT 44.170 -41.550 44.730 -41.380 ;
        RECT 44.170 -43.780 44.340 -41.550 ;
        RECT 44.960 -43.780 45.130 -37.150 ;
        RECT 38.080 -44.340 38.600 -44.170 ;
        RECT 44.570 -44.240 44.740 -43.910 ;
        RECT 38.430 -44.670 38.600 -44.340 ;
        RECT 45.560 -44.700 45.730 -36.700 ;
        RECT 46.000 -44.700 46.170 -36.700 ;
        RECT 46.520 -44.700 46.690 -36.460 ;
        RECT 46.960 -44.700 47.130 -36.700 ;
        RECT 47.490 -44.700 47.660 -36.700 ;
        RECT 47.930 -44.700 48.100 -36.120 ;
        RECT 58.340 -36.290 58.510 -36.060 ;
        RECT 58.690 -36.060 61.450 -35.950 ;
        RECT 68.600 -35.890 68.770 -31.710 ;
        RECT 69.040 -33.660 69.210 -31.710 ;
        RECT 69.040 -33.830 69.250 -33.660 ;
        RECT 69.040 -35.280 69.210 -33.830 ;
        RECT 69.040 -35.450 69.250 -35.280 ;
        RECT 69.040 -35.710 69.210 -35.450 ;
        RECT 70.160 -35.890 70.330 -31.710 ;
        RECT 70.600 -33.650 70.770 -31.710 ;
        RECT 71.130 -33.650 71.300 -31.710 ;
        RECT 70.600 -33.820 71.300 -33.650 ;
        RECT 70.600 -35.270 70.770 -33.820 ;
        RECT 71.130 -35.270 71.300 -33.820 ;
        RECT 70.600 -35.440 70.790 -35.270 ;
        RECT 71.110 -35.440 71.300 -35.270 ;
        RECT 70.600 -35.710 70.770 -35.440 ;
        RECT 71.130 -35.710 71.300 -35.440 ;
        RECT 68.600 -36.060 70.330 -35.890 ;
        RECT 71.570 -35.890 71.740 -31.710 ;
        RECT 72.660 -33.630 72.830 -31.710 ;
        RECT 72.620 -33.800 72.830 -33.630 ;
        RECT 72.660 -35.280 72.830 -33.800 ;
        RECT 72.620 -35.450 72.830 -35.280 ;
        RECT 72.660 -35.710 72.830 -35.450 ;
        RECT 73.100 -35.890 73.270 -31.710 ;
        RECT 73.750 -33.930 73.920 -33.520 ;
        RECT 71.570 -35.950 73.270 -35.890 ;
        RECT 58.690 -36.120 59.920 -36.060 ;
        RECT 48.680 -36.490 49.010 -36.320 ;
        RECT 57.430 -36.500 57.760 -36.330 ;
        RECT 58.340 -36.460 59.580 -36.290 ;
        RECT 48.450 -44.700 48.620 -36.700 ;
        RECT 48.890 -44.700 49.060 -36.700 ;
        RECT 49.850 -36.980 50.020 -36.650 ;
        RECT 56.390 -36.970 56.560 -36.640 ;
        RECT 49.460 -41.140 49.630 -37.150 ;
        RECT 49.900 -37.700 50.070 -37.150 ;
        RECT 56.340 -37.700 56.510 -37.150 ;
        RECT 50.250 -41.140 50.420 -39.140 ;
        RECT 55.990 -41.160 56.160 -39.160 ;
        RECT 49.900 -44.170 50.070 -41.280 ;
        RECT 55.990 -41.550 56.550 -41.380 ;
        RECT 55.990 -43.780 56.160 -41.550 ;
        RECT 56.780 -43.780 56.950 -37.150 ;
        RECT 49.900 -44.340 50.420 -44.170 ;
        RECT 56.390 -44.240 56.560 -43.910 ;
        RECT 50.250 -44.670 50.420 -44.340 ;
        RECT 57.380 -44.700 57.550 -36.700 ;
        RECT 57.820 -44.700 57.990 -36.700 ;
        RECT 58.340 -44.700 58.510 -36.460 ;
        RECT 58.780 -44.700 58.950 -36.700 ;
        RECT 59.310 -44.700 59.480 -36.700 ;
        RECT 59.750 -44.700 59.920 -36.120 ;
        RECT 70.160 -36.290 70.330 -36.060 ;
        RECT 70.510 -36.060 73.270 -35.950 ;
        RECT 80.420 -35.890 80.590 -31.710 ;
        RECT 80.860 -33.660 81.030 -31.710 ;
        RECT 80.860 -33.830 81.070 -33.660 ;
        RECT 80.860 -35.280 81.030 -33.830 ;
        RECT 80.860 -35.450 81.070 -35.280 ;
        RECT 80.860 -35.710 81.030 -35.450 ;
        RECT 81.980 -35.890 82.150 -31.710 ;
        RECT 82.420 -33.650 82.590 -31.710 ;
        RECT 82.950 -33.650 83.120 -31.710 ;
        RECT 82.420 -33.820 83.120 -33.650 ;
        RECT 82.420 -35.270 82.590 -33.820 ;
        RECT 82.950 -35.270 83.120 -33.820 ;
        RECT 82.420 -35.440 82.610 -35.270 ;
        RECT 82.930 -35.440 83.120 -35.270 ;
        RECT 82.420 -35.710 82.590 -35.440 ;
        RECT 82.950 -35.710 83.120 -35.440 ;
        RECT 80.420 -36.060 82.150 -35.890 ;
        RECT 83.390 -35.890 83.560 -31.710 ;
        RECT 84.480 -33.630 84.650 -31.710 ;
        RECT 84.440 -33.800 84.650 -33.630 ;
        RECT 84.480 -35.280 84.650 -33.800 ;
        RECT 84.440 -35.450 84.650 -35.280 ;
        RECT 84.480 -35.710 84.650 -35.450 ;
        RECT 84.920 -35.890 85.090 -31.710 ;
        RECT 85.570 -33.930 85.740 -33.520 ;
        RECT 83.390 -35.950 85.090 -35.890 ;
        RECT 70.510 -36.120 71.740 -36.060 ;
        RECT 60.500 -36.490 60.830 -36.320 ;
        RECT 69.250 -36.500 69.580 -36.330 ;
        RECT 70.160 -36.460 71.400 -36.290 ;
        RECT 60.270 -44.700 60.440 -36.700 ;
        RECT 60.710 -44.700 60.880 -36.700 ;
        RECT 61.670 -36.980 61.840 -36.650 ;
        RECT 68.210 -36.970 68.380 -36.640 ;
        RECT 61.280 -41.140 61.450 -37.150 ;
        RECT 61.720 -37.700 61.890 -37.150 ;
        RECT 68.160 -37.700 68.330 -37.150 ;
        RECT 62.070 -41.140 62.240 -39.140 ;
        RECT 67.810 -41.160 67.980 -39.160 ;
        RECT 61.720 -44.170 61.890 -41.280 ;
        RECT 67.810 -41.550 68.370 -41.380 ;
        RECT 67.810 -43.780 67.980 -41.550 ;
        RECT 68.600 -43.780 68.770 -37.150 ;
        RECT 61.720 -44.340 62.240 -44.170 ;
        RECT 68.210 -44.240 68.380 -43.910 ;
        RECT 62.070 -44.670 62.240 -44.340 ;
        RECT 69.200 -44.700 69.370 -36.700 ;
        RECT 69.640 -44.700 69.810 -36.700 ;
        RECT 70.160 -44.700 70.330 -36.460 ;
        RECT 70.600 -44.700 70.770 -36.700 ;
        RECT 71.130 -44.700 71.300 -36.700 ;
        RECT 71.570 -44.700 71.740 -36.120 ;
        RECT 81.980 -36.290 82.150 -36.060 ;
        RECT 82.330 -36.060 85.090 -35.950 ;
        RECT 92.260 -35.890 92.430 -31.710 ;
        RECT 92.700 -33.660 92.870 -31.710 ;
        RECT 92.700 -33.830 92.910 -33.660 ;
        RECT 92.700 -35.280 92.870 -33.830 ;
        RECT 92.700 -35.450 92.910 -35.280 ;
        RECT 92.700 -35.710 92.870 -35.450 ;
        RECT 93.820 -35.890 93.990 -31.710 ;
        RECT 94.260 -33.650 94.430 -31.710 ;
        RECT 94.790 -33.650 94.960 -31.710 ;
        RECT 94.260 -33.820 94.960 -33.650 ;
        RECT 94.260 -35.270 94.430 -33.820 ;
        RECT 94.790 -35.270 94.960 -33.820 ;
        RECT 94.260 -35.440 94.450 -35.270 ;
        RECT 94.770 -35.440 94.960 -35.270 ;
        RECT 94.260 -35.710 94.430 -35.440 ;
        RECT 94.790 -35.710 94.960 -35.440 ;
        RECT 92.260 -36.060 93.990 -35.890 ;
        RECT 95.230 -35.890 95.400 -31.710 ;
        RECT 96.320 -33.630 96.490 -31.710 ;
        RECT 96.280 -33.800 96.490 -33.630 ;
        RECT 96.320 -35.280 96.490 -33.800 ;
        RECT 96.280 -35.450 96.490 -35.280 ;
        RECT 96.320 -35.710 96.490 -35.450 ;
        RECT 96.760 -35.890 96.930 -31.710 ;
        RECT 97.410 -33.930 97.580 -33.520 ;
        RECT 95.230 -35.950 96.930 -35.890 ;
        RECT 82.330 -36.120 83.560 -36.060 ;
        RECT 72.320 -36.490 72.650 -36.320 ;
        RECT 81.070 -36.500 81.400 -36.330 ;
        RECT 81.980 -36.460 83.220 -36.290 ;
        RECT 72.090 -44.700 72.260 -36.700 ;
        RECT 72.530 -44.700 72.700 -36.700 ;
        RECT 73.490 -36.980 73.660 -36.650 ;
        RECT 80.030 -36.970 80.200 -36.640 ;
        RECT 73.100 -41.140 73.270 -37.150 ;
        RECT 73.540 -37.700 73.710 -37.150 ;
        RECT 79.980 -37.700 80.150 -37.150 ;
        RECT 73.890 -41.140 74.060 -39.140 ;
        RECT 79.630 -41.160 79.800 -39.160 ;
        RECT 73.540 -44.170 73.710 -41.280 ;
        RECT 79.630 -41.550 80.190 -41.380 ;
        RECT 79.630 -43.780 79.800 -41.550 ;
        RECT 80.420 -43.780 80.590 -37.150 ;
        RECT 73.540 -44.340 74.060 -44.170 ;
        RECT 80.030 -44.240 80.200 -43.910 ;
        RECT 73.890 -44.670 74.060 -44.340 ;
        RECT 81.020 -44.700 81.190 -36.700 ;
        RECT 81.460 -44.700 81.630 -36.700 ;
        RECT 81.980 -44.700 82.150 -36.460 ;
        RECT 82.420 -44.700 82.590 -36.700 ;
        RECT 82.950 -44.700 83.120 -36.700 ;
        RECT 83.390 -44.700 83.560 -36.120 ;
        RECT 93.820 -36.290 93.990 -36.060 ;
        RECT 94.170 -36.060 96.930 -35.950 ;
        RECT 104.100 -35.890 104.270 -31.710 ;
        RECT 104.540 -33.660 104.710 -31.710 ;
        RECT 104.540 -33.830 104.750 -33.660 ;
        RECT 104.540 -35.280 104.710 -33.830 ;
        RECT 104.540 -35.450 104.750 -35.280 ;
        RECT 104.540 -35.710 104.710 -35.450 ;
        RECT 105.660 -35.890 105.830 -31.710 ;
        RECT 106.100 -33.650 106.270 -31.710 ;
        RECT 106.630 -33.650 106.800 -31.710 ;
        RECT 106.100 -33.820 106.800 -33.650 ;
        RECT 106.100 -35.270 106.270 -33.820 ;
        RECT 106.630 -35.270 106.800 -33.820 ;
        RECT 106.100 -35.440 106.290 -35.270 ;
        RECT 106.610 -35.440 106.800 -35.270 ;
        RECT 106.100 -35.710 106.270 -35.440 ;
        RECT 106.630 -35.710 106.800 -35.440 ;
        RECT 104.100 -36.060 105.830 -35.890 ;
        RECT 107.070 -35.890 107.240 -31.710 ;
        RECT 108.160 -33.630 108.330 -31.710 ;
        RECT 108.120 -33.800 108.330 -33.630 ;
        RECT 108.160 -35.280 108.330 -33.800 ;
        RECT 108.120 -35.450 108.330 -35.280 ;
        RECT 108.160 -35.710 108.330 -35.450 ;
        RECT 108.600 -35.890 108.770 -31.710 ;
        RECT 109.250 -33.930 109.420 -33.520 ;
        RECT 107.070 -35.950 108.770 -35.890 ;
        RECT 94.170 -36.120 95.400 -36.060 ;
        RECT 84.140 -36.490 84.470 -36.320 ;
        RECT 92.910 -36.500 93.240 -36.330 ;
        RECT 93.820 -36.460 95.060 -36.290 ;
        RECT 83.910 -44.700 84.080 -36.700 ;
        RECT 84.350 -44.700 84.520 -36.700 ;
        RECT 85.310 -36.980 85.480 -36.650 ;
        RECT 91.870 -36.970 92.040 -36.640 ;
        RECT 84.920 -41.140 85.090 -37.150 ;
        RECT 85.360 -37.700 85.530 -37.150 ;
        RECT 91.820 -37.700 91.990 -37.150 ;
        RECT 85.710 -41.140 85.880 -39.140 ;
        RECT 91.470 -41.160 91.640 -39.160 ;
        RECT 85.360 -44.170 85.530 -41.280 ;
        RECT 91.470 -41.550 92.030 -41.380 ;
        RECT 91.470 -43.780 91.640 -41.550 ;
        RECT 92.260 -43.780 92.430 -37.150 ;
        RECT 85.360 -44.340 85.880 -44.170 ;
        RECT 91.870 -44.240 92.040 -43.910 ;
        RECT 85.710 -44.670 85.880 -44.340 ;
        RECT 92.860 -44.700 93.030 -36.700 ;
        RECT 93.300 -44.700 93.470 -36.700 ;
        RECT 93.820 -44.700 93.990 -36.460 ;
        RECT 94.260 -44.700 94.430 -36.700 ;
        RECT 94.790 -44.700 94.960 -36.700 ;
        RECT 95.230 -44.700 95.400 -36.120 ;
        RECT 105.660 -36.290 105.830 -36.060 ;
        RECT 106.010 -36.060 108.770 -35.950 ;
        RECT 115.970 -35.890 116.140 -31.710 ;
        RECT 116.410 -33.660 116.580 -31.710 ;
        RECT 116.410 -33.830 116.620 -33.660 ;
        RECT 116.410 -35.280 116.580 -33.830 ;
        RECT 116.410 -35.450 116.620 -35.280 ;
        RECT 116.410 -35.710 116.580 -35.450 ;
        RECT 117.530 -35.890 117.700 -31.710 ;
        RECT 117.970 -33.650 118.140 -31.710 ;
        RECT 118.500 -33.650 118.670 -31.710 ;
        RECT 117.970 -33.820 118.670 -33.650 ;
        RECT 117.970 -35.270 118.140 -33.820 ;
        RECT 118.500 -35.270 118.670 -33.820 ;
        RECT 117.970 -35.440 118.160 -35.270 ;
        RECT 118.480 -35.440 118.670 -35.270 ;
        RECT 117.970 -35.710 118.140 -35.440 ;
        RECT 118.500 -35.710 118.670 -35.440 ;
        RECT 115.970 -36.060 117.700 -35.890 ;
        RECT 118.940 -35.890 119.110 -31.710 ;
        RECT 120.030 -33.630 120.200 -31.710 ;
        RECT 119.990 -33.800 120.200 -33.630 ;
        RECT 120.030 -35.280 120.200 -33.800 ;
        RECT 119.990 -35.450 120.200 -35.280 ;
        RECT 120.030 -35.710 120.200 -35.450 ;
        RECT 120.470 -35.890 120.640 -31.710 ;
        RECT 121.120 -33.930 121.290 -33.520 ;
        RECT 118.940 -35.950 120.640 -35.890 ;
        RECT 106.010 -36.120 107.240 -36.060 ;
        RECT 95.980 -36.490 96.310 -36.320 ;
        RECT 104.750 -36.500 105.080 -36.330 ;
        RECT 105.660 -36.460 106.900 -36.290 ;
        RECT 95.750 -44.700 95.920 -36.700 ;
        RECT 96.190 -44.700 96.360 -36.700 ;
        RECT 97.150 -36.980 97.320 -36.650 ;
        RECT 103.710 -36.970 103.880 -36.640 ;
        RECT 96.760 -41.140 96.930 -37.150 ;
        RECT 97.200 -37.700 97.370 -37.150 ;
        RECT 103.660 -37.700 103.830 -37.150 ;
        RECT 97.550 -41.140 97.720 -39.140 ;
        RECT 103.310 -41.160 103.480 -39.160 ;
        RECT 97.200 -44.170 97.370 -41.280 ;
        RECT 103.310 -41.550 103.870 -41.380 ;
        RECT 103.310 -43.780 103.480 -41.550 ;
        RECT 104.100 -43.780 104.270 -37.150 ;
        RECT 97.200 -44.340 97.720 -44.170 ;
        RECT 103.710 -44.240 103.880 -43.910 ;
        RECT 97.550 -44.670 97.720 -44.340 ;
        RECT 104.700 -44.700 104.870 -36.700 ;
        RECT 105.140 -44.700 105.310 -36.700 ;
        RECT 105.660 -44.700 105.830 -36.460 ;
        RECT 106.100 -44.700 106.270 -36.700 ;
        RECT 106.630 -44.700 106.800 -36.700 ;
        RECT 107.070 -44.700 107.240 -36.120 ;
        RECT 117.530 -36.290 117.700 -36.060 ;
        RECT 117.880 -36.060 120.640 -35.950 ;
        RECT 127.840 -35.890 128.010 -31.710 ;
        RECT 128.280 -33.660 128.450 -31.710 ;
        RECT 128.280 -33.830 128.490 -33.660 ;
        RECT 128.280 -35.280 128.450 -33.830 ;
        RECT 128.280 -35.450 128.490 -35.280 ;
        RECT 128.280 -35.710 128.450 -35.450 ;
        RECT 129.400 -35.890 129.570 -31.710 ;
        RECT 129.840 -33.650 130.010 -31.710 ;
        RECT 130.370 -33.650 130.540 -31.710 ;
        RECT 129.840 -33.820 130.540 -33.650 ;
        RECT 129.840 -35.270 130.010 -33.820 ;
        RECT 130.370 -35.270 130.540 -33.820 ;
        RECT 129.840 -35.440 130.030 -35.270 ;
        RECT 130.350 -35.440 130.540 -35.270 ;
        RECT 129.840 -35.710 130.010 -35.440 ;
        RECT 130.370 -35.710 130.540 -35.440 ;
        RECT 127.840 -36.060 129.570 -35.890 ;
        RECT 130.810 -35.890 130.980 -31.710 ;
        RECT 131.900 -33.630 132.070 -31.710 ;
        RECT 131.860 -33.800 132.070 -33.630 ;
        RECT 131.900 -35.280 132.070 -33.800 ;
        RECT 131.860 -35.450 132.070 -35.280 ;
        RECT 131.900 -35.710 132.070 -35.450 ;
        RECT 132.340 -35.890 132.510 -31.710 ;
        RECT 132.990 -33.930 133.160 -33.520 ;
        RECT 130.810 -35.950 132.510 -35.890 ;
        RECT 117.880 -36.120 119.110 -36.060 ;
        RECT 107.820 -36.490 108.150 -36.320 ;
        RECT 116.620 -36.500 116.950 -36.330 ;
        RECT 117.530 -36.460 118.770 -36.290 ;
        RECT 107.590 -44.700 107.760 -36.700 ;
        RECT 108.030 -44.700 108.200 -36.700 ;
        RECT 108.990 -36.980 109.160 -36.650 ;
        RECT 115.580 -36.970 115.750 -36.640 ;
        RECT 108.600 -41.140 108.770 -37.150 ;
        RECT 109.040 -37.700 109.210 -37.150 ;
        RECT 115.530 -37.700 115.700 -37.150 ;
        RECT 109.390 -41.140 109.560 -39.140 ;
        RECT 115.180 -41.160 115.350 -39.160 ;
        RECT 109.040 -44.170 109.210 -41.280 ;
        RECT 115.180 -41.550 115.740 -41.380 ;
        RECT 115.180 -43.780 115.350 -41.550 ;
        RECT 115.970 -43.780 116.140 -37.150 ;
        RECT 109.040 -44.340 109.560 -44.170 ;
        RECT 115.580 -44.240 115.750 -43.910 ;
        RECT 109.390 -44.670 109.560 -44.340 ;
        RECT 116.570 -44.700 116.740 -36.700 ;
        RECT 117.010 -44.700 117.180 -36.700 ;
        RECT 117.530 -44.700 117.700 -36.460 ;
        RECT 117.970 -44.700 118.140 -36.700 ;
        RECT 118.500 -44.700 118.670 -36.700 ;
        RECT 118.940 -44.700 119.110 -36.120 ;
        RECT 129.400 -36.290 129.570 -36.060 ;
        RECT 129.750 -36.060 132.510 -35.950 ;
        RECT 136.850 -35.890 137.020 -31.710 ;
        RECT 137.290 -33.660 137.460 -31.710 ;
        RECT 137.290 -33.830 137.500 -33.660 ;
        RECT 137.290 -35.280 137.460 -33.830 ;
        RECT 137.290 -35.450 137.500 -35.280 ;
        RECT 137.290 -35.710 137.460 -35.450 ;
        RECT 138.410 -35.890 138.580 -31.710 ;
        RECT 138.850 -33.650 139.020 -31.710 ;
        RECT 139.380 -33.650 139.550 -31.710 ;
        RECT 138.850 -33.820 139.550 -33.650 ;
        RECT 138.850 -35.270 139.020 -33.820 ;
        RECT 139.380 -35.270 139.550 -33.820 ;
        RECT 138.850 -35.440 139.040 -35.270 ;
        RECT 139.360 -35.440 139.550 -35.270 ;
        RECT 138.850 -35.710 139.020 -35.440 ;
        RECT 139.380 -35.710 139.550 -35.440 ;
        RECT 136.850 -36.060 138.580 -35.890 ;
        RECT 139.820 -35.890 139.990 -31.710 ;
        RECT 140.910 -33.630 141.080 -31.710 ;
        RECT 140.870 -33.800 141.080 -33.630 ;
        RECT 140.910 -35.280 141.080 -33.800 ;
        RECT 140.870 -35.450 141.080 -35.280 ;
        RECT 140.910 -35.710 141.080 -35.450 ;
        RECT 141.350 -35.890 141.520 -31.710 ;
        RECT 142.000 -33.930 142.170 -33.520 ;
        RECT 139.820 -35.950 141.520 -35.890 ;
        RECT 129.750 -36.120 130.980 -36.060 ;
        RECT 119.690 -36.490 120.020 -36.320 ;
        RECT 128.490 -36.500 128.820 -36.330 ;
        RECT 129.400 -36.460 130.640 -36.290 ;
        RECT 119.460 -44.700 119.630 -36.700 ;
        RECT 119.900 -44.700 120.070 -36.700 ;
        RECT 120.860 -36.980 121.030 -36.650 ;
        RECT 127.450 -36.970 127.620 -36.640 ;
        RECT 120.470 -41.140 120.640 -37.150 ;
        RECT 120.910 -37.700 121.080 -37.150 ;
        RECT 127.400 -37.700 127.570 -37.150 ;
        RECT 121.260 -41.140 121.430 -39.140 ;
        RECT 127.050 -41.160 127.220 -39.160 ;
        RECT 120.910 -44.170 121.080 -41.280 ;
        RECT 127.050 -41.550 127.610 -41.380 ;
        RECT 127.050 -43.780 127.220 -41.550 ;
        RECT 127.840 -43.780 128.010 -37.150 ;
        RECT 120.910 -44.340 121.430 -44.170 ;
        RECT 127.450 -44.240 127.620 -43.910 ;
        RECT 121.260 -44.670 121.430 -44.340 ;
        RECT 128.440 -44.700 128.610 -36.700 ;
        RECT 128.880 -44.700 129.050 -36.700 ;
        RECT 129.400 -44.700 129.570 -36.460 ;
        RECT 129.840 -44.700 130.010 -36.700 ;
        RECT 130.370 -44.700 130.540 -36.700 ;
        RECT 130.810 -44.700 130.980 -36.120 ;
        RECT 138.410 -36.290 138.580 -36.060 ;
        RECT 138.760 -36.060 141.520 -35.950 ;
        RECT 138.760 -36.120 139.990 -36.060 ;
        RECT 131.560 -36.490 131.890 -36.320 ;
        RECT 137.500 -36.500 137.830 -36.330 ;
        RECT 138.410 -36.460 139.650 -36.290 ;
        RECT 131.330 -44.700 131.500 -36.700 ;
        RECT 131.770 -44.700 131.940 -36.700 ;
        RECT 132.730 -36.980 132.900 -36.650 ;
        RECT 136.460 -36.970 136.630 -36.640 ;
        RECT 132.340 -41.140 132.510 -37.150 ;
        RECT 132.780 -37.700 132.950 -37.150 ;
        RECT 136.410 -37.700 136.580 -37.150 ;
        RECT 133.130 -41.140 133.300 -39.140 ;
        RECT 136.060 -41.160 136.230 -39.160 ;
        RECT 132.780 -44.170 132.950 -41.280 ;
        RECT 136.060 -41.550 136.620 -41.380 ;
        RECT 136.060 -43.780 136.230 -41.550 ;
        RECT 136.850 -43.780 137.020 -37.150 ;
        RECT 132.780 -44.340 133.300 -44.170 ;
        RECT 136.460 -44.240 136.630 -43.910 ;
        RECT 133.130 -44.670 133.300 -44.340 ;
        RECT 137.450 -44.700 137.620 -36.700 ;
        RECT 137.890 -44.700 138.060 -36.700 ;
        RECT 138.410 -44.700 138.580 -36.460 ;
        RECT 138.850 -44.700 139.020 -36.700 ;
        RECT 139.380 -44.700 139.550 -36.700 ;
        RECT 139.820 -44.700 139.990 -36.120 ;
        RECT 140.570 -36.490 140.900 -36.320 ;
        RECT 140.340 -44.700 140.510 -36.700 ;
        RECT 140.780 -44.700 140.950 -36.700 ;
        RECT 141.740 -36.980 141.910 -36.650 ;
        RECT 141.350 -41.140 141.520 -37.150 ;
        RECT 141.790 -37.700 141.960 -37.150 ;
        RECT 142.140 -41.140 142.310 -39.140 ;
        RECT 141.790 -44.170 141.960 -41.280 ;
        RECT 141.790 -44.340 142.310 -44.170 ;
        RECT 142.140 -44.670 142.310 -44.340 ;
        RECT -32.820 -45.300 -32.650 -44.890 ;
        RECT -21.320 -45.300 -21.150 -44.890 ;
        RECT -9.500 -45.300 -9.330 -44.890 ;
        RECT 2.310 -45.300 2.480 -44.890 ;
        RECT 14.120 -45.300 14.290 -44.890 ;
        RECT 25.940 -45.300 26.110 -44.890 ;
        RECT 37.760 -45.300 37.930 -44.890 ;
        RECT 49.580 -45.300 49.750 -44.890 ;
        RECT 61.400 -45.300 61.570 -44.890 ;
        RECT 73.220 -45.300 73.390 -44.890 ;
        RECT 85.040 -45.300 85.210 -44.890 ;
        RECT 96.880 -45.300 97.050 -44.890 ;
        RECT 108.720 -45.300 108.890 -44.890 ;
        RECT 120.590 -45.300 120.760 -44.890 ;
        RECT 132.460 -45.300 132.630 -44.890 ;
        RECT 141.470 -45.300 141.640 -44.890 ;
        RECT -37.830 -48.790 -37.660 -48.460 ;
        RECT -38.230 -50.920 -38.060 -48.920 ;
        RECT -37.880 -52.930 -37.710 -52.380 ;
        RECT -37.440 -52.930 -37.270 -46.380 ;
        RECT -37.830 -53.440 -37.660 -53.110 ;
        RECT -36.840 -53.380 -36.670 -45.380 ;
        RECT -36.400 -53.380 -36.230 -45.380 ;
        RECT -36.790 -53.750 -36.460 -53.580 ;
        RECT -35.880 -53.620 -35.710 -45.380 ;
        RECT -35.440 -53.380 -35.270 -45.380 ;
        RECT -34.910 -53.380 -34.740 -45.380 ;
        RECT -35.880 -53.790 -34.640 -53.620 ;
        RECT -36.320 -54.020 -36.150 -54.010 ;
        RECT -35.880 -54.020 -35.710 -53.790 ;
        RECT -34.470 -53.960 -34.300 -45.380 ;
        RECT -33.950 -53.380 -33.780 -45.380 ;
        RECT -33.510 -53.380 -33.340 -45.380 ;
        RECT -32.150 -45.720 -31.980 -45.400 ;
        RECT -32.500 -45.890 -31.980 -45.720 ;
        RECT -32.500 -48.820 -32.330 -45.890 ;
        RECT -26.330 -48.790 -26.160 -48.460 ;
        RECT -32.940 -52.930 -32.770 -48.940 ;
        RECT -32.150 -50.940 -31.980 -48.940 ;
        RECT -26.730 -50.920 -26.560 -48.920 ;
        RECT -32.500 -52.930 -32.330 -52.380 ;
        RECT -26.380 -52.930 -26.210 -52.380 ;
        RECT -25.940 -52.930 -25.770 -46.380 ;
        RECT -32.550 -53.430 -32.380 -53.100 ;
        RECT -26.330 -53.440 -26.160 -53.110 ;
        RECT -25.340 -53.380 -25.170 -45.380 ;
        RECT -24.900 -53.380 -24.730 -45.380 ;
        RECT -33.720 -53.760 -33.390 -53.590 ;
        RECT -25.290 -53.750 -24.960 -53.580 ;
        RECT -24.380 -53.620 -24.210 -45.380 ;
        RECT -23.940 -53.380 -23.770 -45.380 ;
        RECT -23.410 -53.380 -23.240 -45.380 ;
        RECT -37.440 -54.190 -35.710 -54.020 ;
        RECT -35.530 -54.020 -34.300 -53.960 ;
        RECT -24.380 -53.790 -23.140 -53.620 ;
        RECT -24.380 -54.020 -24.210 -53.790 ;
        RECT -22.970 -53.960 -22.800 -45.380 ;
        RECT -22.450 -53.380 -22.280 -45.380 ;
        RECT -22.010 -53.380 -21.840 -45.380 ;
        RECT -20.650 -45.720 -20.480 -45.390 ;
        RECT -21.000 -45.890 -20.480 -45.720 ;
        RECT -21.000 -48.820 -20.830 -45.890 ;
        RECT -14.510 -48.790 -14.340 -48.460 ;
        RECT -21.440 -52.930 -21.270 -48.940 ;
        RECT -20.650 -50.940 -20.480 -48.940 ;
        RECT -14.910 -50.920 -14.740 -48.920 ;
        RECT -21.000 -52.930 -20.830 -52.380 ;
        RECT -14.560 -52.930 -14.390 -52.380 ;
        RECT -14.120 -52.930 -13.950 -46.380 ;
        RECT -21.050 -53.430 -20.880 -53.100 ;
        RECT -14.510 -53.440 -14.340 -53.110 ;
        RECT -13.520 -53.380 -13.350 -45.380 ;
        RECT -13.080 -53.380 -12.910 -45.380 ;
        RECT -22.220 -53.760 -21.890 -53.590 ;
        RECT -13.470 -53.750 -13.140 -53.580 ;
        RECT -12.560 -53.620 -12.390 -45.380 ;
        RECT -12.120 -53.380 -11.950 -45.380 ;
        RECT -11.590 -53.380 -11.420 -45.380 ;
        RECT -35.530 -54.130 -32.770 -54.020 ;
        RECT -37.440 -58.370 -37.270 -54.190 ;
        RECT -37.000 -54.630 -36.830 -54.370 ;
        RECT -37.000 -54.800 -36.790 -54.630 ;
        RECT -37.000 -56.250 -36.830 -54.800 ;
        RECT -37.000 -56.420 -36.790 -56.250 ;
        RECT -37.000 -58.370 -36.830 -56.420 ;
        RECT -35.880 -58.370 -35.710 -54.190 ;
        RECT -34.470 -54.190 -32.770 -54.130 ;
        RECT -35.440 -54.640 -35.270 -54.370 ;
        RECT -34.910 -54.640 -34.740 -54.370 ;
        RECT -35.440 -54.810 -35.250 -54.640 ;
        RECT -34.930 -54.810 -34.740 -54.640 ;
        RECT -35.440 -56.260 -35.270 -54.810 ;
        RECT -34.910 -56.260 -34.740 -54.810 ;
        RECT -35.440 -56.430 -34.740 -56.260 ;
        RECT -35.440 -58.370 -35.270 -56.430 ;
        RECT -34.910 -58.370 -34.740 -56.430 ;
        RECT -34.470 -58.370 -34.300 -54.190 ;
        RECT -33.380 -54.630 -33.210 -54.370 ;
        RECT -33.420 -54.800 -33.210 -54.630 ;
        RECT -33.380 -56.280 -33.210 -54.800 ;
        RECT -33.420 -56.450 -33.210 -56.280 ;
        RECT -33.380 -58.370 -33.210 -56.450 ;
        RECT -32.940 -58.370 -32.770 -54.190 ;
        RECT -25.940 -54.190 -24.210 -54.020 ;
        RECT -24.030 -54.020 -22.800 -53.960 ;
        RECT -12.560 -53.790 -11.320 -53.620 ;
        RECT -12.560 -54.020 -12.390 -53.790 ;
        RECT -11.150 -53.960 -10.980 -45.380 ;
        RECT -10.630 -53.380 -10.460 -45.380 ;
        RECT -10.190 -53.380 -10.020 -45.380 ;
        RECT -8.830 -45.720 -8.660 -45.390 ;
        RECT -9.180 -45.890 -8.660 -45.720 ;
        RECT -9.180 -48.820 -9.010 -45.890 ;
        RECT -2.700 -48.790 -2.530 -48.460 ;
        RECT -9.620 -52.930 -9.450 -48.940 ;
        RECT -8.830 -50.940 -8.660 -48.940 ;
        RECT -3.100 -50.920 -2.930 -48.920 ;
        RECT -9.180 -52.930 -9.010 -52.380 ;
        RECT -2.750 -52.930 -2.580 -52.380 ;
        RECT -2.310 -52.930 -2.140 -46.380 ;
        RECT -9.230 -53.430 -9.060 -53.100 ;
        RECT -2.700 -53.440 -2.530 -53.110 ;
        RECT -1.710 -53.380 -1.540 -45.380 ;
        RECT -1.270 -53.380 -1.100 -45.380 ;
        RECT -10.400 -53.760 -10.070 -53.590 ;
        RECT -1.660 -53.750 -1.330 -53.580 ;
        RECT -0.750 -53.620 -0.580 -45.380 ;
        RECT -0.310 -53.380 -0.140 -45.380 ;
        RECT 0.220 -53.380 0.390 -45.380 ;
        RECT -24.030 -54.130 -21.270 -54.020 ;
        RECT -32.290 -56.550 -32.120 -56.140 ;
        RECT -25.940 -58.370 -25.770 -54.190 ;
        RECT -25.500 -54.630 -25.330 -54.370 ;
        RECT -25.500 -54.800 -25.290 -54.630 ;
        RECT -25.500 -56.250 -25.330 -54.800 ;
        RECT -25.500 -56.420 -25.290 -56.250 ;
        RECT -25.500 -58.370 -25.330 -56.420 ;
        RECT -24.380 -58.370 -24.210 -54.190 ;
        RECT -22.970 -54.190 -21.270 -54.130 ;
        RECT -23.940 -54.640 -23.770 -54.370 ;
        RECT -23.410 -54.640 -23.240 -54.370 ;
        RECT -23.940 -54.810 -23.750 -54.640 ;
        RECT -23.430 -54.810 -23.240 -54.640 ;
        RECT -23.940 -56.260 -23.770 -54.810 ;
        RECT -23.410 -56.260 -23.240 -54.810 ;
        RECT -23.940 -56.430 -23.240 -56.260 ;
        RECT -23.940 -58.370 -23.770 -56.430 ;
        RECT -23.410 -58.370 -23.240 -56.430 ;
        RECT -22.970 -58.370 -22.800 -54.190 ;
        RECT -21.880 -54.630 -21.710 -54.370 ;
        RECT -21.920 -54.800 -21.710 -54.630 ;
        RECT -21.880 -56.280 -21.710 -54.800 ;
        RECT -21.920 -56.450 -21.710 -56.280 ;
        RECT -21.880 -58.370 -21.710 -56.450 ;
        RECT -21.440 -58.370 -21.270 -54.190 ;
        RECT -14.120 -54.190 -12.390 -54.020 ;
        RECT -12.210 -54.020 -10.980 -53.960 ;
        RECT -0.750 -53.790 0.490 -53.620 ;
        RECT -0.750 -54.020 -0.580 -53.790 ;
        RECT 0.660 -53.960 0.830 -45.380 ;
        RECT 1.180 -53.380 1.350 -45.380 ;
        RECT 1.620 -53.380 1.790 -45.380 ;
        RECT 2.980 -45.720 3.150 -45.390 ;
        RECT 2.630 -45.890 3.150 -45.720 ;
        RECT 2.630 -48.820 2.800 -45.890 ;
        RECT 9.110 -48.790 9.280 -48.460 ;
        RECT 2.190 -52.930 2.360 -48.940 ;
        RECT 2.980 -50.940 3.150 -48.940 ;
        RECT 8.710 -50.920 8.880 -48.920 ;
        RECT 2.630 -52.930 2.800 -52.380 ;
        RECT 9.060 -52.930 9.230 -52.380 ;
        RECT 9.500 -52.930 9.670 -46.380 ;
        RECT 2.580 -53.430 2.750 -53.100 ;
        RECT 9.110 -53.440 9.280 -53.110 ;
        RECT 10.100 -53.380 10.270 -45.380 ;
        RECT 10.540 -53.380 10.710 -45.380 ;
        RECT 1.410 -53.760 1.740 -53.590 ;
        RECT 10.150 -53.750 10.480 -53.580 ;
        RECT 11.060 -53.620 11.230 -45.380 ;
        RECT 11.500 -53.380 11.670 -45.380 ;
        RECT 12.030 -53.380 12.200 -45.380 ;
        RECT -12.210 -54.130 -9.450 -54.020 ;
        RECT -20.790 -56.550 -20.620 -56.140 ;
        RECT -14.120 -58.370 -13.950 -54.190 ;
        RECT -13.680 -54.630 -13.510 -54.370 ;
        RECT -13.680 -54.800 -13.470 -54.630 ;
        RECT -13.680 -56.250 -13.510 -54.800 ;
        RECT -13.680 -56.420 -13.470 -56.250 ;
        RECT -13.680 -58.370 -13.510 -56.420 ;
        RECT -12.560 -58.370 -12.390 -54.190 ;
        RECT -11.150 -54.190 -9.450 -54.130 ;
        RECT -12.120 -54.640 -11.950 -54.370 ;
        RECT -11.590 -54.640 -11.420 -54.370 ;
        RECT -12.120 -54.810 -11.930 -54.640 ;
        RECT -11.610 -54.810 -11.420 -54.640 ;
        RECT -12.120 -56.260 -11.950 -54.810 ;
        RECT -11.590 -56.260 -11.420 -54.810 ;
        RECT -12.120 -56.430 -11.420 -56.260 ;
        RECT -12.120 -58.370 -11.950 -56.430 ;
        RECT -11.590 -58.370 -11.420 -56.430 ;
        RECT -11.150 -58.370 -10.980 -54.190 ;
        RECT -10.060 -54.630 -9.890 -54.370 ;
        RECT -10.100 -54.800 -9.890 -54.630 ;
        RECT -10.060 -56.280 -9.890 -54.800 ;
        RECT -10.100 -56.450 -9.890 -56.280 ;
        RECT -10.060 -58.370 -9.890 -56.450 ;
        RECT -9.620 -58.370 -9.450 -54.190 ;
        RECT -2.310 -54.190 -0.580 -54.020 ;
        RECT -0.400 -54.020 0.830 -53.960 ;
        RECT 11.060 -53.790 12.300 -53.620 ;
        RECT 11.060 -54.020 11.230 -53.790 ;
        RECT 12.470 -53.960 12.640 -45.380 ;
        RECT 12.990 -53.380 13.160 -45.380 ;
        RECT 13.430 -53.380 13.600 -45.380 ;
        RECT 14.790 -45.720 14.960 -45.390 ;
        RECT 14.440 -45.890 14.960 -45.720 ;
        RECT 14.440 -48.820 14.610 -45.890 ;
        RECT 20.930 -48.790 21.100 -48.460 ;
        RECT 14.000 -52.930 14.170 -48.940 ;
        RECT 14.790 -50.940 14.960 -48.940 ;
        RECT 20.530 -50.920 20.700 -48.920 ;
        RECT 14.440 -52.930 14.610 -52.380 ;
        RECT 20.880 -52.930 21.050 -52.380 ;
        RECT 21.320 -52.930 21.490 -46.380 ;
        RECT 14.390 -53.430 14.560 -53.100 ;
        RECT 20.930 -53.440 21.100 -53.110 ;
        RECT 21.920 -53.380 22.090 -45.380 ;
        RECT 22.360 -53.380 22.530 -45.380 ;
        RECT 13.220 -53.760 13.550 -53.590 ;
        RECT 21.970 -53.750 22.300 -53.580 ;
        RECT 22.880 -53.620 23.050 -45.380 ;
        RECT 23.320 -53.380 23.490 -45.380 ;
        RECT 23.850 -53.380 24.020 -45.380 ;
        RECT -0.400 -54.130 2.360 -54.020 ;
        RECT -8.970 -56.550 -8.800 -56.140 ;
        RECT -2.310 -58.370 -2.140 -54.190 ;
        RECT -1.870 -54.630 -1.700 -54.370 ;
        RECT -1.870 -54.800 -1.660 -54.630 ;
        RECT -1.870 -56.250 -1.700 -54.800 ;
        RECT -1.870 -56.420 -1.660 -56.250 ;
        RECT -1.870 -58.370 -1.700 -56.420 ;
        RECT -0.750 -58.370 -0.580 -54.190 ;
        RECT 0.660 -54.190 2.360 -54.130 ;
        RECT -0.310 -54.640 -0.140 -54.370 ;
        RECT 0.220 -54.640 0.390 -54.370 ;
        RECT -0.310 -54.810 -0.120 -54.640 ;
        RECT 0.200 -54.810 0.390 -54.640 ;
        RECT -0.310 -56.260 -0.140 -54.810 ;
        RECT 0.220 -56.260 0.390 -54.810 ;
        RECT -0.310 -56.430 0.390 -56.260 ;
        RECT -0.310 -58.370 -0.140 -56.430 ;
        RECT 0.220 -58.370 0.390 -56.430 ;
        RECT 0.660 -58.370 0.830 -54.190 ;
        RECT 1.750 -54.630 1.920 -54.370 ;
        RECT 1.710 -54.800 1.920 -54.630 ;
        RECT 1.750 -56.280 1.920 -54.800 ;
        RECT 1.710 -56.450 1.920 -56.280 ;
        RECT 1.750 -58.370 1.920 -56.450 ;
        RECT 2.190 -58.370 2.360 -54.190 ;
        RECT 9.500 -54.190 11.230 -54.020 ;
        RECT 11.410 -54.020 12.640 -53.960 ;
        RECT 22.880 -53.790 24.120 -53.620 ;
        RECT 22.880 -54.020 23.050 -53.790 ;
        RECT 24.290 -53.960 24.460 -45.380 ;
        RECT 24.810 -53.380 24.980 -45.380 ;
        RECT 25.250 -53.380 25.420 -45.380 ;
        RECT 26.610 -45.720 26.780 -45.390 ;
        RECT 26.260 -45.890 26.780 -45.720 ;
        RECT 26.260 -48.820 26.430 -45.890 ;
        RECT 32.750 -48.790 32.920 -48.460 ;
        RECT 25.820 -52.930 25.990 -48.940 ;
        RECT 26.610 -50.940 26.780 -48.940 ;
        RECT 32.350 -50.920 32.520 -48.920 ;
        RECT 26.260 -52.930 26.430 -52.380 ;
        RECT 32.700 -52.930 32.870 -52.380 ;
        RECT 33.140 -52.930 33.310 -46.380 ;
        RECT 26.210 -53.430 26.380 -53.100 ;
        RECT 32.750 -53.440 32.920 -53.110 ;
        RECT 33.740 -53.380 33.910 -45.380 ;
        RECT 34.180 -53.380 34.350 -45.380 ;
        RECT 25.040 -53.760 25.370 -53.590 ;
        RECT 33.790 -53.750 34.120 -53.580 ;
        RECT 34.700 -53.620 34.870 -45.380 ;
        RECT 35.140 -53.380 35.310 -45.380 ;
        RECT 35.670 -53.380 35.840 -45.380 ;
        RECT 11.410 -54.130 14.170 -54.020 ;
        RECT 2.840 -56.550 3.010 -56.140 ;
        RECT 9.500 -58.370 9.670 -54.190 ;
        RECT 9.940 -54.630 10.110 -54.370 ;
        RECT 9.940 -54.800 10.150 -54.630 ;
        RECT 9.940 -56.250 10.110 -54.800 ;
        RECT 9.940 -56.420 10.150 -56.250 ;
        RECT 9.940 -58.370 10.110 -56.420 ;
        RECT 11.060 -58.370 11.230 -54.190 ;
        RECT 12.470 -54.190 14.170 -54.130 ;
        RECT 11.500 -54.640 11.670 -54.370 ;
        RECT 12.030 -54.640 12.200 -54.370 ;
        RECT 11.500 -54.810 11.690 -54.640 ;
        RECT 12.010 -54.810 12.200 -54.640 ;
        RECT 11.500 -56.260 11.670 -54.810 ;
        RECT 12.030 -56.260 12.200 -54.810 ;
        RECT 11.500 -56.430 12.200 -56.260 ;
        RECT 11.500 -58.370 11.670 -56.430 ;
        RECT 12.030 -58.370 12.200 -56.430 ;
        RECT 12.470 -58.370 12.640 -54.190 ;
        RECT 13.560 -54.630 13.730 -54.370 ;
        RECT 13.520 -54.800 13.730 -54.630 ;
        RECT 13.560 -56.280 13.730 -54.800 ;
        RECT 13.520 -56.450 13.730 -56.280 ;
        RECT 13.560 -58.370 13.730 -56.450 ;
        RECT 14.000 -58.370 14.170 -54.190 ;
        RECT 21.320 -54.190 23.050 -54.020 ;
        RECT 23.230 -54.020 24.460 -53.960 ;
        RECT 34.700 -53.790 35.940 -53.620 ;
        RECT 34.700 -54.020 34.870 -53.790 ;
        RECT 36.110 -53.960 36.280 -45.380 ;
        RECT 36.630 -53.380 36.800 -45.380 ;
        RECT 37.070 -53.380 37.240 -45.380 ;
        RECT 38.430 -45.720 38.600 -45.390 ;
        RECT 38.080 -45.890 38.600 -45.720 ;
        RECT 38.080 -48.820 38.250 -45.890 ;
        RECT 44.570 -48.790 44.740 -48.460 ;
        RECT 37.640 -52.930 37.810 -48.940 ;
        RECT 38.430 -50.940 38.600 -48.940 ;
        RECT 44.170 -50.920 44.340 -48.920 ;
        RECT 38.080 -52.930 38.250 -52.380 ;
        RECT 44.520 -52.930 44.690 -52.380 ;
        RECT 44.960 -52.930 45.130 -46.380 ;
        RECT 38.030 -53.430 38.200 -53.100 ;
        RECT 44.570 -53.440 44.740 -53.110 ;
        RECT 45.560 -53.380 45.730 -45.380 ;
        RECT 46.000 -53.380 46.170 -45.380 ;
        RECT 36.860 -53.760 37.190 -53.590 ;
        RECT 45.610 -53.750 45.940 -53.580 ;
        RECT 46.520 -53.620 46.690 -45.380 ;
        RECT 46.960 -53.380 47.130 -45.380 ;
        RECT 47.490 -53.380 47.660 -45.380 ;
        RECT 23.230 -54.130 25.990 -54.020 ;
        RECT 14.650 -56.550 14.820 -56.140 ;
        RECT 21.320 -58.370 21.490 -54.190 ;
        RECT 21.760 -54.630 21.930 -54.370 ;
        RECT 21.760 -54.800 21.970 -54.630 ;
        RECT 21.760 -56.250 21.930 -54.800 ;
        RECT 21.760 -56.420 21.970 -56.250 ;
        RECT 21.760 -58.370 21.930 -56.420 ;
        RECT 22.880 -58.370 23.050 -54.190 ;
        RECT 24.290 -54.190 25.990 -54.130 ;
        RECT 23.320 -54.640 23.490 -54.370 ;
        RECT 23.850 -54.640 24.020 -54.370 ;
        RECT 23.320 -54.810 23.510 -54.640 ;
        RECT 23.830 -54.810 24.020 -54.640 ;
        RECT 23.320 -56.260 23.490 -54.810 ;
        RECT 23.850 -56.260 24.020 -54.810 ;
        RECT 23.320 -56.430 24.020 -56.260 ;
        RECT 23.320 -58.370 23.490 -56.430 ;
        RECT 23.850 -58.370 24.020 -56.430 ;
        RECT 24.290 -58.370 24.460 -54.190 ;
        RECT 25.380 -54.630 25.550 -54.370 ;
        RECT 25.340 -54.800 25.550 -54.630 ;
        RECT 25.380 -56.280 25.550 -54.800 ;
        RECT 25.340 -56.450 25.550 -56.280 ;
        RECT 25.380 -58.370 25.550 -56.450 ;
        RECT 25.820 -58.370 25.990 -54.190 ;
        RECT 33.140 -54.190 34.870 -54.020 ;
        RECT 35.050 -54.020 36.280 -53.960 ;
        RECT 46.520 -53.790 47.760 -53.620 ;
        RECT 46.520 -54.020 46.690 -53.790 ;
        RECT 47.930 -53.960 48.100 -45.380 ;
        RECT 48.450 -53.380 48.620 -45.380 ;
        RECT 48.890 -53.380 49.060 -45.380 ;
        RECT 50.250 -45.720 50.420 -45.390 ;
        RECT 49.900 -45.890 50.420 -45.720 ;
        RECT 49.900 -48.820 50.070 -45.890 ;
        RECT 56.390 -48.790 56.560 -48.460 ;
        RECT 49.460 -52.930 49.630 -48.940 ;
        RECT 50.250 -50.940 50.420 -48.940 ;
        RECT 55.990 -50.920 56.160 -48.920 ;
        RECT 49.900 -52.930 50.070 -52.380 ;
        RECT 56.340 -52.930 56.510 -52.380 ;
        RECT 56.780 -52.930 56.950 -46.380 ;
        RECT 49.850 -53.430 50.020 -53.100 ;
        RECT 56.390 -53.440 56.560 -53.110 ;
        RECT 57.380 -53.380 57.550 -45.380 ;
        RECT 57.820 -53.380 57.990 -45.380 ;
        RECT 48.680 -53.760 49.010 -53.590 ;
        RECT 57.430 -53.750 57.760 -53.580 ;
        RECT 58.340 -53.620 58.510 -45.380 ;
        RECT 58.780 -53.380 58.950 -45.380 ;
        RECT 59.310 -53.380 59.480 -45.380 ;
        RECT 35.050 -54.130 37.810 -54.020 ;
        RECT 26.470 -56.550 26.640 -56.140 ;
        RECT 33.140 -58.370 33.310 -54.190 ;
        RECT 33.580 -54.630 33.750 -54.370 ;
        RECT 33.580 -54.800 33.790 -54.630 ;
        RECT 33.580 -56.250 33.750 -54.800 ;
        RECT 33.580 -56.420 33.790 -56.250 ;
        RECT 33.580 -58.370 33.750 -56.420 ;
        RECT 34.700 -58.370 34.870 -54.190 ;
        RECT 36.110 -54.190 37.810 -54.130 ;
        RECT 35.140 -54.640 35.310 -54.370 ;
        RECT 35.670 -54.640 35.840 -54.370 ;
        RECT 35.140 -54.810 35.330 -54.640 ;
        RECT 35.650 -54.810 35.840 -54.640 ;
        RECT 35.140 -56.260 35.310 -54.810 ;
        RECT 35.670 -56.260 35.840 -54.810 ;
        RECT 35.140 -56.430 35.840 -56.260 ;
        RECT 35.140 -58.370 35.310 -56.430 ;
        RECT 35.670 -58.370 35.840 -56.430 ;
        RECT 36.110 -58.370 36.280 -54.190 ;
        RECT 37.200 -54.630 37.370 -54.370 ;
        RECT 37.160 -54.800 37.370 -54.630 ;
        RECT 37.200 -56.280 37.370 -54.800 ;
        RECT 37.160 -56.450 37.370 -56.280 ;
        RECT 37.200 -58.370 37.370 -56.450 ;
        RECT 37.640 -58.370 37.810 -54.190 ;
        RECT 44.960 -54.190 46.690 -54.020 ;
        RECT 46.870 -54.020 48.100 -53.960 ;
        RECT 58.340 -53.790 59.580 -53.620 ;
        RECT 58.340 -54.020 58.510 -53.790 ;
        RECT 59.750 -53.960 59.920 -45.380 ;
        RECT 60.270 -53.380 60.440 -45.380 ;
        RECT 60.710 -53.380 60.880 -45.380 ;
        RECT 62.070 -45.720 62.240 -45.390 ;
        RECT 61.720 -45.890 62.240 -45.720 ;
        RECT 61.720 -48.820 61.890 -45.890 ;
        RECT 68.210 -48.790 68.380 -48.460 ;
        RECT 61.280 -52.930 61.450 -48.940 ;
        RECT 62.070 -50.940 62.240 -48.940 ;
        RECT 67.810 -50.920 67.980 -48.920 ;
        RECT 61.720 -52.930 61.890 -52.380 ;
        RECT 68.160 -52.930 68.330 -52.380 ;
        RECT 68.600 -52.930 68.770 -46.380 ;
        RECT 61.670 -53.430 61.840 -53.100 ;
        RECT 68.210 -53.440 68.380 -53.110 ;
        RECT 69.200 -53.380 69.370 -45.380 ;
        RECT 69.640 -53.380 69.810 -45.380 ;
        RECT 60.500 -53.760 60.830 -53.590 ;
        RECT 69.250 -53.750 69.580 -53.580 ;
        RECT 70.160 -53.620 70.330 -45.380 ;
        RECT 70.600 -53.380 70.770 -45.380 ;
        RECT 71.130 -53.380 71.300 -45.380 ;
        RECT 46.870 -54.130 49.630 -54.020 ;
        RECT 38.290 -56.550 38.460 -56.140 ;
        RECT 44.960 -58.370 45.130 -54.190 ;
        RECT 45.400 -54.630 45.570 -54.370 ;
        RECT 45.400 -54.800 45.610 -54.630 ;
        RECT 45.400 -56.250 45.570 -54.800 ;
        RECT 45.400 -56.420 45.610 -56.250 ;
        RECT 45.400 -58.370 45.570 -56.420 ;
        RECT 46.520 -58.370 46.690 -54.190 ;
        RECT 47.930 -54.190 49.630 -54.130 ;
        RECT 46.960 -54.640 47.130 -54.370 ;
        RECT 47.490 -54.640 47.660 -54.370 ;
        RECT 46.960 -54.810 47.150 -54.640 ;
        RECT 47.470 -54.810 47.660 -54.640 ;
        RECT 46.960 -56.260 47.130 -54.810 ;
        RECT 47.490 -56.260 47.660 -54.810 ;
        RECT 46.960 -56.430 47.660 -56.260 ;
        RECT 46.960 -58.370 47.130 -56.430 ;
        RECT 47.490 -58.370 47.660 -56.430 ;
        RECT 47.930 -58.370 48.100 -54.190 ;
        RECT 49.020 -54.630 49.190 -54.370 ;
        RECT 48.980 -54.800 49.190 -54.630 ;
        RECT 49.020 -56.280 49.190 -54.800 ;
        RECT 48.980 -56.450 49.190 -56.280 ;
        RECT 49.020 -58.370 49.190 -56.450 ;
        RECT 49.460 -58.370 49.630 -54.190 ;
        RECT 56.780 -54.190 58.510 -54.020 ;
        RECT 58.690 -54.020 59.920 -53.960 ;
        RECT 70.160 -53.790 71.400 -53.620 ;
        RECT 70.160 -54.020 70.330 -53.790 ;
        RECT 71.570 -53.960 71.740 -45.380 ;
        RECT 72.090 -53.380 72.260 -45.380 ;
        RECT 72.530 -53.380 72.700 -45.380 ;
        RECT 73.890 -45.720 74.060 -45.390 ;
        RECT 73.540 -45.890 74.060 -45.720 ;
        RECT 73.540 -48.820 73.710 -45.890 ;
        RECT 80.030 -48.790 80.200 -48.460 ;
        RECT 73.100 -52.930 73.270 -48.940 ;
        RECT 73.890 -50.940 74.060 -48.940 ;
        RECT 79.630 -50.920 79.800 -48.920 ;
        RECT 73.540 -52.930 73.710 -52.380 ;
        RECT 79.980 -52.930 80.150 -52.380 ;
        RECT 80.420 -52.930 80.590 -46.380 ;
        RECT 73.490 -53.430 73.660 -53.100 ;
        RECT 80.030 -53.440 80.200 -53.110 ;
        RECT 81.020 -53.380 81.190 -45.380 ;
        RECT 81.460 -53.380 81.630 -45.380 ;
        RECT 72.320 -53.760 72.650 -53.590 ;
        RECT 81.070 -53.750 81.400 -53.580 ;
        RECT 81.980 -53.620 82.150 -45.380 ;
        RECT 82.420 -53.380 82.590 -45.380 ;
        RECT 82.950 -53.380 83.120 -45.380 ;
        RECT 58.690 -54.130 61.450 -54.020 ;
        RECT 50.110 -56.550 50.280 -56.140 ;
        RECT 56.780 -58.370 56.950 -54.190 ;
        RECT 57.220 -54.630 57.390 -54.370 ;
        RECT 57.220 -54.800 57.430 -54.630 ;
        RECT 57.220 -56.250 57.390 -54.800 ;
        RECT 57.220 -56.420 57.430 -56.250 ;
        RECT 57.220 -58.370 57.390 -56.420 ;
        RECT 58.340 -58.370 58.510 -54.190 ;
        RECT 59.750 -54.190 61.450 -54.130 ;
        RECT 58.780 -54.640 58.950 -54.370 ;
        RECT 59.310 -54.640 59.480 -54.370 ;
        RECT 58.780 -54.810 58.970 -54.640 ;
        RECT 59.290 -54.810 59.480 -54.640 ;
        RECT 58.780 -56.260 58.950 -54.810 ;
        RECT 59.310 -56.260 59.480 -54.810 ;
        RECT 58.780 -56.430 59.480 -56.260 ;
        RECT 58.780 -58.370 58.950 -56.430 ;
        RECT 59.310 -58.370 59.480 -56.430 ;
        RECT 59.750 -58.370 59.920 -54.190 ;
        RECT 60.840 -54.630 61.010 -54.370 ;
        RECT 60.800 -54.800 61.010 -54.630 ;
        RECT 60.840 -56.280 61.010 -54.800 ;
        RECT 60.800 -56.450 61.010 -56.280 ;
        RECT 60.840 -58.370 61.010 -56.450 ;
        RECT 61.280 -58.370 61.450 -54.190 ;
        RECT 68.600 -54.190 70.330 -54.020 ;
        RECT 70.510 -54.020 71.740 -53.960 ;
        RECT 81.980 -53.790 83.220 -53.620 ;
        RECT 81.980 -54.020 82.150 -53.790 ;
        RECT 83.390 -53.960 83.560 -45.380 ;
        RECT 83.910 -53.380 84.080 -45.380 ;
        RECT 84.350 -53.380 84.520 -45.380 ;
        RECT 85.710 -45.720 85.880 -45.390 ;
        RECT 85.360 -45.890 85.880 -45.720 ;
        RECT 85.360 -48.820 85.530 -45.890 ;
        RECT 91.870 -48.790 92.040 -48.460 ;
        RECT 84.920 -52.930 85.090 -48.940 ;
        RECT 85.710 -50.940 85.880 -48.940 ;
        RECT 91.470 -50.920 91.640 -48.920 ;
        RECT 85.360 -52.930 85.530 -52.380 ;
        RECT 91.820 -52.930 91.990 -52.380 ;
        RECT 92.260 -52.930 92.430 -46.380 ;
        RECT 85.310 -53.430 85.480 -53.100 ;
        RECT 91.870 -53.440 92.040 -53.110 ;
        RECT 92.860 -53.380 93.030 -45.380 ;
        RECT 93.300 -53.380 93.470 -45.380 ;
        RECT 84.140 -53.760 84.470 -53.590 ;
        RECT 92.910 -53.750 93.240 -53.580 ;
        RECT 93.820 -53.620 93.990 -45.380 ;
        RECT 94.260 -53.380 94.430 -45.380 ;
        RECT 94.790 -53.380 94.960 -45.380 ;
        RECT 70.510 -54.130 73.270 -54.020 ;
        RECT 61.930 -56.550 62.100 -56.140 ;
        RECT 68.600 -58.370 68.770 -54.190 ;
        RECT 69.040 -54.630 69.210 -54.370 ;
        RECT 69.040 -54.800 69.250 -54.630 ;
        RECT 69.040 -56.250 69.210 -54.800 ;
        RECT 69.040 -56.420 69.250 -56.250 ;
        RECT 69.040 -58.370 69.210 -56.420 ;
        RECT 70.160 -58.370 70.330 -54.190 ;
        RECT 71.570 -54.190 73.270 -54.130 ;
        RECT 70.600 -54.640 70.770 -54.370 ;
        RECT 71.130 -54.640 71.300 -54.370 ;
        RECT 70.600 -54.810 70.790 -54.640 ;
        RECT 71.110 -54.810 71.300 -54.640 ;
        RECT 70.600 -56.260 70.770 -54.810 ;
        RECT 71.130 -56.260 71.300 -54.810 ;
        RECT 70.600 -56.430 71.300 -56.260 ;
        RECT 70.600 -58.370 70.770 -56.430 ;
        RECT 71.130 -58.370 71.300 -56.430 ;
        RECT 71.570 -58.370 71.740 -54.190 ;
        RECT 72.660 -54.630 72.830 -54.370 ;
        RECT 72.620 -54.800 72.830 -54.630 ;
        RECT 72.660 -56.280 72.830 -54.800 ;
        RECT 72.620 -56.450 72.830 -56.280 ;
        RECT 72.660 -58.370 72.830 -56.450 ;
        RECT 73.100 -58.370 73.270 -54.190 ;
        RECT 80.420 -54.190 82.150 -54.020 ;
        RECT 82.330 -54.020 83.560 -53.960 ;
        RECT 93.820 -53.790 95.060 -53.620 ;
        RECT 93.820 -54.020 93.990 -53.790 ;
        RECT 95.230 -53.960 95.400 -45.380 ;
        RECT 95.750 -53.380 95.920 -45.380 ;
        RECT 96.190 -53.380 96.360 -45.380 ;
        RECT 97.550 -45.720 97.720 -45.390 ;
        RECT 97.200 -45.890 97.720 -45.720 ;
        RECT 97.200 -48.820 97.370 -45.890 ;
        RECT 103.710 -48.790 103.880 -48.460 ;
        RECT 96.760 -52.930 96.930 -48.940 ;
        RECT 97.550 -50.940 97.720 -48.940 ;
        RECT 103.310 -50.920 103.480 -48.920 ;
        RECT 97.200 -52.930 97.370 -52.380 ;
        RECT 103.660 -52.930 103.830 -52.380 ;
        RECT 104.100 -52.930 104.270 -46.380 ;
        RECT 97.150 -53.430 97.320 -53.100 ;
        RECT 103.710 -53.440 103.880 -53.110 ;
        RECT 104.700 -53.380 104.870 -45.380 ;
        RECT 105.140 -53.380 105.310 -45.380 ;
        RECT 95.980 -53.760 96.310 -53.590 ;
        RECT 104.750 -53.750 105.080 -53.580 ;
        RECT 105.660 -53.620 105.830 -45.380 ;
        RECT 106.100 -53.380 106.270 -45.380 ;
        RECT 106.630 -53.380 106.800 -45.380 ;
        RECT 82.330 -54.130 85.090 -54.020 ;
        RECT 73.750 -56.550 73.920 -56.140 ;
        RECT 80.420 -58.370 80.590 -54.190 ;
        RECT 80.860 -54.630 81.030 -54.370 ;
        RECT 80.860 -54.800 81.070 -54.630 ;
        RECT 80.860 -56.250 81.030 -54.800 ;
        RECT 80.860 -56.420 81.070 -56.250 ;
        RECT 80.860 -58.370 81.030 -56.420 ;
        RECT 81.980 -58.370 82.150 -54.190 ;
        RECT 83.390 -54.190 85.090 -54.130 ;
        RECT 82.420 -54.640 82.590 -54.370 ;
        RECT 82.950 -54.640 83.120 -54.370 ;
        RECT 82.420 -54.810 82.610 -54.640 ;
        RECT 82.930 -54.810 83.120 -54.640 ;
        RECT 82.420 -56.260 82.590 -54.810 ;
        RECT 82.950 -56.260 83.120 -54.810 ;
        RECT 82.420 -56.430 83.120 -56.260 ;
        RECT 82.420 -58.370 82.590 -56.430 ;
        RECT 82.950 -58.370 83.120 -56.430 ;
        RECT 83.390 -58.370 83.560 -54.190 ;
        RECT 84.480 -54.630 84.650 -54.370 ;
        RECT 84.440 -54.800 84.650 -54.630 ;
        RECT 84.480 -56.280 84.650 -54.800 ;
        RECT 84.440 -56.450 84.650 -56.280 ;
        RECT 84.480 -58.370 84.650 -56.450 ;
        RECT 84.920 -58.370 85.090 -54.190 ;
        RECT 92.260 -54.190 93.990 -54.020 ;
        RECT 94.170 -54.020 95.400 -53.960 ;
        RECT 105.660 -53.790 106.900 -53.620 ;
        RECT 105.660 -54.020 105.830 -53.790 ;
        RECT 107.070 -53.960 107.240 -45.380 ;
        RECT 107.590 -53.380 107.760 -45.380 ;
        RECT 108.030 -53.380 108.200 -45.380 ;
        RECT 109.390 -45.720 109.560 -45.400 ;
        RECT 109.040 -45.890 109.560 -45.720 ;
        RECT 109.040 -48.820 109.210 -45.890 ;
        RECT 115.580 -48.790 115.750 -48.460 ;
        RECT 108.600 -52.930 108.770 -48.940 ;
        RECT 109.390 -50.940 109.560 -48.940 ;
        RECT 115.180 -50.920 115.350 -48.920 ;
        RECT 109.040 -52.930 109.210 -52.380 ;
        RECT 115.530 -52.930 115.700 -52.380 ;
        RECT 115.970 -52.930 116.140 -46.380 ;
        RECT 108.990 -53.430 109.160 -53.100 ;
        RECT 115.580 -53.440 115.750 -53.110 ;
        RECT 116.570 -53.380 116.740 -45.380 ;
        RECT 117.010 -53.380 117.180 -45.380 ;
        RECT 107.820 -53.760 108.150 -53.590 ;
        RECT 116.620 -53.750 116.950 -53.580 ;
        RECT 117.530 -53.620 117.700 -45.380 ;
        RECT 117.970 -53.380 118.140 -45.380 ;
        RECT 118.500 -53.380 118.670 -45.380 ;
        RECT 94.170 -54.130 96.930 -54.020 ;
        RECT 85.570 -56.550 85.740 -56.140 ;
        RECT 92.260 -58.370 92.430 -54.190 ;
        RECT 92.700 -54.630 92.870 -54.370 ;
        RECT 92.700 -54.800 92.910 -54.630 ;
        RECT 92.700 -56.250 92.870 -54.800 ;
        RECT 92.700 -56.420 92.910 -56.250 ;
        RECT 92.700 -58.370 92.870 -56.420 ;
        RECT 93.820 -58.370 93.990 -54.190 ;
        RECT 95.230 -54.190 96.930 -54.130 ;
        RECT 94.260 -54.640 94.430 -54.370 ;
        RECT 94.790 -54.640 94.960 -54.370 ;
        RECT 94.260 -54.810 94.450 -54.640 ;
        RECT 94.770 -54.810 94.960 -54.640 ;
        RECT 94.260 -56.260 94.430 -54.810 ;
        RECT 94.790 -56.260 94.960 -54.810 ;
        RECT 94.260 -56.430 94.960 -56.260 ;
        RECT 94.260 -58.370 94.430 -56.430 ;
        RECT 94.790 -58.370 94.960 -56.430 ;
        RECT 95.230 -58.370 95.400 -54.190 ;
        RECT 96.320 -54.630 96.490 -54.370 ;
        RECT 96.280 -54.800 96.490 -54.630 ;
        RECT 96.320 -56.280 96.490 -54.800 ;
        RECT 96.280 -56.450 96.490 -56.280 ;
        RECT 96.320 -58.370 96.490 -56.450 ;
        RECT 96.760 -58.370 96.930 -54.190 ;
        RECT 104.100 -54.190 105.830 -54.020 ;
        RECT 106.010 -54.020 107.240 -53.960 ;
        RECT 117.530 -53.790 118.770 -53.620 ;
        RECT 117.530 -54.020 117.700 -53.790 ;
        RECT 118.940 -53.960 119.110 -45.380 ;
        RECT 119.460 -53.380 119.630 -45.380 ;
        RECT 119.900 -53.380 120.070 -45.380 ;
        RECT 121.260 -45.720 121.430 -45.390 ;
        RECT 120.910 -45.890 121.430 -45.720 ;
        RECT 120.910 -48.820 121.080 -45.890 ;
        RECT 127.450 -48.790 127.620 -48.460 ;
        RECT 120.470 -52.930 120.640 -48.940 ;
        RECT 121.260 -50.940 121.430 -48.940 ;
        RECT 127.050 -50.920 127.220 -48.920 ;
        RECT 120.910 -52.930 121.080 -52.380 ;
        RECT 127.400 -52.930 127.570 -52.380 ;
        RECT 127.840 -52.930 128.010 -46.380 ;
        RECT 120.860 -53.430 121.030 -53.100 ;
        RECT 127.450 -53.440 127.620 -53.110 ;
        RECT 128.440 -53.380 128.610 -45.380 ;
        RECT 128.880 -53.380 129.050 -45.380 ;
        RECT 119.690 -53.760 120.020 -53.590 ;
        RECT 128.490 -53.750 128.820 -53.580 ;
        RECT 129.400 -53.620 129.570 -45.380 ;
        RECT 129.840 -53.380 130.010 -45.380 ;
        RECT 130.370 -53.380 130.540 -45.380 ;
        RECT 106.010 -54.130 108.770 -54.020 ;
        RECT 97.410 -56.550 97.580 -56.140 ;
        RECT 104.100 -58.370 104.270 -54.190 ;
        RECT 104.540 -54.630 104.710 -54.370 ;
        RECT 104.540 -54.800 104.750 -54.630 ;
        RECT 104.540 -56.250 104.710 -54.800 ;
        RECT 104.540 -56.420 104.750 -56.250 ;
        RECT 104.540 -58.370 104.710 -56.420 ;
        RECT 105.660 -58.370 105.830 -54.190 ;
        RECT 107.070 -54.190 108.770 -54.130 ;
        RECT 106.100 -54.640 106.270 -54.370 ;
        RECT 106.630 -54.640 106.800 -54.370 ;
        RECT 106.100 -54.810 106.290 -54.640 ;
        RECT 106.610 -54.810 106.800 -54.640 ;
        RECT 106.100 -56.260 106.270 -54.810 ;
        RECT 106.630 -56.260 106.800 -54.810 ;
        RECT 106.100 -56.430 106.800 -56.260 ;
        RECT 106.100 -58.370 106.270 -56.430 ;
        RECT 106.630 -58.370 106.800 -56.430 ;
        RECT 107.070 -58.370 107.240 -54.190 ;
        RECT 108.160 -54.630 108.330 -54.370 ;
        RECT 108.120 -54.800 108.330 -54.630 ;
        RECT 108.160 -56.280 108.330 -54.800 ;
        RECT 108.120 -56.450 108.330 -56.280 ;
        RECT 108.160 -58.370 108.330 -56.450 ;
        RECT 108.600 -58.370 108.770 -54.190 ;
        RECT 115.970 -54.190 117.700 -54.020 ;
        RECT 117.880 -54.020 119.110 -53.960 ;
        RECT 129.400 -53.790 130.640 -53.620 ;
        RECT 129.400 -54.020 129.570 -53.790 ;
        RECT 130.810 -53.960 130.980 -45.380 ;
        RECT 131.330 -53.380 131.500 -45.380 ;
        RECT 131.770 -53.380 131.940 -45.380 ;
        RECT 133.130 -45.720 133.300 -45.390 ;
        RECT 132.780 -45.890 133.300 -45.720 ;
        RECT 132.780 -48.820 132.950 -45.890 ;
        RECT 136.460 -48.790 136.630 -48.460 ;
        RECT 132.340 -52.930 132.510 -48.940 ;
        RECT 133.130 -50.940 133.300 -48.940 ;
        RECT 136.060 -50.920 136.230 -48.920 ;
        RECT 132.780 -52.930 132.950 -52.380 ;
        RECT 136.410 -52.930 136.580 -52.380 ;
        RECT 136.850 -52.930 137.020 -46.380 ;
        RECT 132.730 -53.430 132.900 -53.100 ;
        RECT 136.460 -53.440 136.630 -53.110 ;
        RECT 137.450 -53.380 137.620 -45.380 ;
        RECT 137.890 -53.380 138.060 -45.380 ;
        RECT 131.560 -53.760 131.890 -53.590 ;
        RECT 137.500 -53.750 137.830 -53.580 ;
        RECT 138.410 -53.620 138.580 -45.380 ;
        RECT 138.850 -53.380 139.020 -45.380 ;
        RECT 139.380 -53.380 139.550 -45.380 ;
        RECT 117.880 -54.130 120.640 -54.020 ;
        RECT 109.250 -56.550 109.420 -56.140 ;
        RECT 115.970 -58.370 116.140 -54.190 ;
        RECT 116.410 -54.630 116.580 -54.370 ;
        RECT 116.410 -54.800 116.620 -54.630 ;
        RECT 116.410 -56.250 116.580 -54.800 ;
        RECT 116.410 -56.420 116.620 -56.250 ;
        RECT 116.410 -58.370 116.580 -56.420 ;
        RECT 117.530 -58.370 117.700 -54.190 ;
        RECT 118.940 -54.190 120.640 -54.130 ;
        RECT 117.970 -54.640 118.140 -54.370 ;
        RECT 118.500 -54.640 118.670 -54.370 ;
        RECT 117.970 -54.810 118.160 -54.640 ;
        RECT 118.480 -54.810 118.670 -54.640 ;
        RECT 117.970 -56.260 118.140 -54.810 ;
        RECT 118.500 -56.260 118.670 -54.810 ;
        RECT 117.970 -56.430 118.670 -56.260 ;
        RECT 117.970 -58.370 118.140 -56.430 ;
        RECT 118.500 -58.370 118.670 -56.430 ;
        RECT 118.940 -58.370 119.110 -54.190 ;
        RECT 120.030 -54.630 120.200 -54.370 ;
        RECT 119.990 -54.800 120.200 -54.630 ;
        RECT 120.030 -56.280 120.200 -54.800 ;
        RECT 119.990 -56.450 120.200 -56.280 ;
        RECT 120.030 -58.370 120.200 -56.450 ;
        RECT 120.470 -58.370 120.640 -54.190 ;
        RECT 127.840 -54.190 129.570 -54.020 ;
        RECT 129.750 -54.020 130.980 -53.960 ;
        RECT 138.410 -53.790 139.650 -53.620 ;
        RECT 138.410 -54.020 138.580 -53.790 ;
        RECT 139.820 -53.960 139.990 -45.380 ;
        RECT 140.340 -53.380 140.510 -45.380 ;
        RECT 140.780 -53.380 140.950 -45.380 ;
        RECT 142.140 -45.720 142.310 -45.390 ;
        RECT 141.790 -45.890 142.310 -45.720 ;
        RECT 141.790 -48.820 141.960 -45.890 ;
        RECT 141.350 -52.930 141.520 -48.940 ;
        RECT 142.140 -50.940 142.310 -48.940 ;
        RECT 141.790 -52.930 141.960 -52.380 ;
        RECT 141.740 -53.430 141.910 -53.100 ;
        RECT 140.570 -53.760 140.900 -53.590 ;
        RECT 129.750 -54.130 132.510 -54.020 ;
        RECT 121.120 -56.550 121.290 -56.140 ;
        RECT 127.840 -58.370 128.010 -54.190 ;
        RECT 128.280 -54.630 128.450 -54.370 ;
        RECT 128.280 -54.800 128.490 -54.630 ;
        RECT 128.280 -56.250 128.450 -54.800 ;
        RECT 128.280 -56.420 128.490 -56.250 ;
        RECT 128.280 -58.370 128.450 -56.420 ;
        RECT 129.400 -58.370 129.570 -54.190 ;
        RECT 130.810 -54.190 132.510 -54.130 ;
        RECT 129.840 -54.640 130.010 -54.370 ;
        RECT 130.370 -54.640 130.540 -54.370 ;
        RECT 129.840 -54.810 130.030 -54.640 ;
        RECT 130.350 -54.810 130.540 -54.640 ;
        RECT 129.840 -56.260 130.010 -54.810 ;
        RECT 130.370 -56.260 130.540 -54.810 ;
        RECT 129.840 -56.430 130.540 -56.260 ;
        RECT 129.840 -58.370 130.010 -56.430 ;
        RECT 130.370 -58.370 130.540 -56.430 ;
        RECT 130.810 -58.370 130.980 -54.190 ;
        RECT 131.900 -54.630 132.070 -54.370 ;
        RECT 131.860 -54.800 132.070 -54.630 ;
        RECT 131.900 -56.280 132.070 -54.800 ;
        RECT 131.860 -56.450 132.070 -56.280 ;
        RECT 131.900 -58.370 132.070 -56.450 ;
        RECT 132.340 -58.370 132.510 -54.190 ;
        RECT 136.850 -54.190 138.580 -54.020 ;
        RECT 138.760 -54.020 139.990 -53.960 ;
        RECT 138.760 -54.130 141.520 -54.020 ;
        RECT 132.990 -56.550 133.160 -56.140 ;
        RECT 136.850 -58.370 137.020 -54.190 ;
        RECT 137.290 -54.630 137.460 -54.370 ;
        RECT 137.290 -54.800 137.500 -54.630 ;
        RECT 137.290 -56.250 137.460 -54.800 ;
        RECT 137.290 -56.420 137.500 -56.250 ;
        RECT 137.290 -58.370 137.460 -56.420 ;
        RECT 138.410 -58.370 138.580 -54.190 ;
        RECT 139.820 -54.190 141.520 -54.130 ;
        RECT 138.850 -54.640 139.020 -54.370 ;
        RECT 139.380 -54.640 139.550 -54.370 ;
        RECT 138.850 -54.810 139.040 -54.640 ;
        RECT 139.360 -54.810 139.550 -54.640 ;
        RECT 138.850 -56.260 139.020 -54.810 ;
        RECT 139.380 -56.260 139.550 -54.810 ;
        RECT 138.850 -56.430 139.550 -56.260 ;
        RECT 138.850 -58.370 139.020 -56.430 ;
        RECT 139.380 -58.370 139.550 -56.430 ;
        RECT 139.820 -58.370 139.990 -54.190 ;
        RECT 140.910 -54.630 141.080 -54.370 ;
        RECT 140.870 -54.800 141.080 -54.630 ;
        RECT 140.910 -56.280 141.080 -54.800 ;
        RECT 140.870 -56.450 141.080 -56.280 ;
        RECT 140.910 -58.370 141.080 -56.450 ;
        RECT 141.350 -58.370 141.520 -54.190 ;
        RECT 142.000 -56.550 142.170 -56.140 ;
        RECT -37.290 -58.790 -36.960 -58.620 ;
        RECT -33.240 -58.790 -32.910 -58.620 ;
        RECT -25.790 -58.790 -25.460 -58.620 ;
        RECT -21.740 -58.790 -21.410 -58.620 ;
        RECT -13.970 -58.790 -13.640 -58.620 ;
        RECT -9.920 -58.790 -9.590 -58.620 ;
        RECT -2.160 -58.790 -1.830 -58.620 ;
        RECT 1.890 -58.790 2.220 -58.620 ;
        RECT 9.650 -58.790 9.980 -58.620 ;
        RECT 13.700 -58.790 14.030 -58.620 ;
        RECT 21.470 -58.790 21.800 -58.620 ;
        RECT 25.520 -58.790 25.850 -58.620 ;
        RECT 33.290 -58.790 33.620 -58.620 ;
        RECT 37.340 -58.790 37.670 -58.620 ;
        RECT 45.110 -58.790 45.440 -58.620 ;
        RECT 49.160 -58.790 49.490 -58.620 ;
        RECT 56.930 -58.790 57.260 -58.620 ;
        RECT 60.980 -58.790 61.310 -58.620 ;
        RECT 68.750 -58.790 69.080 -58.620 ;
        RECT 72.800 -58.790 73.130 -58.620 ;
        RECT 80.570 -58.790 80.900 -58.620 ;
        RECT 84.620 -58.790 84.950 -58.620 ;
        RECT 92.410 -58.790 92.740 -58.620 ;
        RECT 96.460 -58.790 96.790 -58.620 ;
        RECT 104.250 -58.790 104.580 -58.620 ;
        RECT 108.300 -58.790 108.630 -58.620 ;
        RECT 116.120 -58.790 116.450 -58.620 ;
        RECT 120.170 -58.790 120.500 -58.620 ;
        RECT 127.990 -58.790 128.320 -58.620 ;
        RECT 132.040 -58.790 132.370 -58.620 ;
        RECT 137.000 -58.790 137.330 -58.620 ;
        RECT 141.050 -58.790 141.380 -58.620 ;
        RECT -37.440 -63.220 -37.270 -59.040 ;
        RECT -37.000 -60.990 -36.830 -59.040 ;
        RECT -37.000 -61.160 -36.790 -60.990 ;
        RECT -37.000 -62.610 -36.830 -61.160 ;
        RECT -37.000 -62.780 -36.790 -62.610 ;
        RECT -37.000 -63.040 -36.830 -62.780 ;
        RECT -35.880 -63.220 -35.710 -59.040 ;
        RECT -35.440 -60.980 -35.270 -59.040 ;
        RECT -34.910 -60.980 -34.740 -59.040 ;
        RECT -35.440 -61.150 -34.740 -60.980 ;
        RECT -35.440 -62.600 -35.270 -61.150 ;
        RECT -34.910 -62.600 -34.740 -61.150 ;
        RECT -35.440 -62.770 -35.250 -62.600 ;
        RECT -34.930 -62.770 -34.740 -62.600 ;
        RECT -35.440 -63.040 -35.270 -62.770 ;
        RECT -34.910 -63.040 -34.740 -62.770 ;
        RECT -37.440 -63.390 -35.710 -63.220 ;
        RECT -34.470 -63.220 -34.300 -59.040 ;
        RECT -33.380 -60.960 -33.210 -59.040 ;
        RECT -33.420 -61.130 -33.210 -60.960 ;
        RECT -33.380 -62.610 -33.210 -61.130 ;
        RECT -33.420 -62.780 -33.210 -62.610 ;
        RECT -33.380 -63.040 -33.210 -62.780 ;
        RECT -32.940 -63.220 -32.770 -59.040 ;
        RECT -32.300 -61.260 -32.130 -60.850 ;
        RECT -34.470 -63.280 -32.770 -63.220 ;
        RECT -35.880 -63.620 -35.710 -63.390 ;
        RECT -35.530 -63.390 -32.770 -63.280 ;
        RECT -25.940 -63.220 -25.770 -59.040 ;
        RECT -25.500 -60.990 -25.330 -59.040 ;
        RECT -25.500 -61.160 -25.290 -60.990 ;
        RECT -25.500 -62.610 -25.330 -61.160 ;
        RECT -25.500 -62.780 -25.290 -62.610 ;
        RECT -25.500 -63.040 -25.330 -62.780 ;
        RECT -24.380 -63.220 -24.210 -59.040 ;
        RECT -23.940 -60.980 -23.770 -59.040 ;
        RECT -23.410 -60.980 -23.240 -59.040 ;
        RECT -23.940 -61.150 -23.240 -60.980 ;
        RECT -23.940 -62.600 -23.770 -61.150 ;
        RECT -23.410 -62.600 -23.240 -61.150 ;
        RECT -23.940 -62.770 -23.750 -62.600 ;
        RECT -23.430 -62.770 -23.240 -62.600 ;
        RECT -23.940 -63.040 -23.770 -62.770 ;
        RECT -23.410 -63.040 -23.240 -62.770 ;
        RECT -25.940 -63.390 -24.210 -63.220 ;
        RECT -22.970 -63.220 -22.800 -59.040 ;
        RECT -21.880 -60.960 -21.710 -59.040 ;
        RECT -21.920 -61.130 -21.710 -60.960 ;
        RECT -21.880 -62.610 -21.710 -61.130 ;
        RECT -21.920 -62.780 -21.710 -62.610 ;
        RECT -21.880 -63.040 -21.710 -62.780 ;
        RECT -21.440 -63.220 -21.270 -59.040 ;
        RECT -20.800 -61.260 -20.630 -60.850 ;
        RECT -22.970 -63.280 -21.270 -63.220 ;
        RECT -35.530 -63.450 -34.300 -63.390 ;
        RECT -36.790 -63.830 -36.460 -63.660 ;
        RECT -35.880 -63.790 -34.640 -63.620 ;
        RECT -37.830 -64.300 -37.660 -63.970 ;
        RECT -37.880 -65.030 -37.710 -64.480 ;
        RECT -37.830 -66.360 -37.660 -66.030 ;
        RECT -38.230 -68.490 -38.060 -66.490 ;
        RECT -37.840 -68.950 -37.670 -68.620 ;
        RECT -37.440 -71.030 -37.270 -64.480 ;
        RECT -36.840 -72.030 -36.670 -64.030 ;
        RECT -36.400 -72.030 -36.230 -64.030 ;
        RECT -35.880 -72.030 -35.710 -63.790 ;
        RECT -35.440 -72.030 -35.270 -64.030 ;
        RECT -34.910 -72.030 -34.740 -64.030 ;
        RECT -34.470 -72.030 -34.300 -63.450 ;
        RECT -24.380 -63.620 -24.210 -63.390 ;
        RECT -24.030 -63.390 -21.270 -63.280 ;
        RECT -14.120 -63.220 -13.950 -59.040 ;
        RECT -13.680 -60.990 -13.510 -59.040 ;
        RECT -13.680 -61.160 -13.470 -60.990 ;
        RECT -13.680 -62.610 -13.510 -61.160 ;
        RECT -13.680 -62.780 -13.470 -62.610 ;
        RECT -13.680 -63.040 -13.510 -62.780 ;
        RECT -12.560 -63.220 -12.390 -59.040 ;
        RECT -12.120 -60.980 -11.950 -59.040 ;
        RECT -11.590 -60.980 -11.420 -59.040 ;
        RECT -12.120 -61.150 -11.420 -60.980 ;
        RECT -12.120 -62.600 -11.950 -61.150 ;
        RECT -11.590 -62.600 -11.420 -61.150 ;
        RECT -12.120 -62.770 -11.930 -62.600 ;
        RECT -11.610 -62.770 -11.420 -62.600 ;
        RECT -12.120 -63.040 -11.950 -62.770 ;
        RECT -11.590 -63.040 -11.420 -62.770 ;
        RECT -14.120 -63.390 -12.390 -63.220 ;
        RECT -11.150 -63.220 -10.980 -59.040 ;
        RECT -10.060 -60.960 -9.890 -59.040 ;
        RECT -10.100 -61.130 -9.890 -60.960 ;
        RECT -10.060 -62.610 -9.890 -61.130 ;
        RECT -10.100 -62.780 -9.890 -62.610 ;
        RECT -10.060 -63.040 -9.890 -62.780 ;
        RECT -9.620 -63.220 -9.450 -59.040 ;
        RECT -8.980 -61.260 -8.810 -60.850 ;
        RECT -11.150 -63.280 -9.450 -63.220 ;
        RECT -24.030 -63.450 -22.800 -63.390 ;
        RECT -33.720 -63.820 -33.390 -63.650 ;
        RECT -25.290 -63.830 -24.960 -63.660 ;
        RECT -24.380 -63.790 -23.140 -63.620 ;
        RECT -33.950 -72.030 -33.780 -64.030 ;
        RECT -33.510 -72.030 -33.340 -64.030 ;
        RECT -32.550 -64.310 -32.380 -63.980 ;
        RECT -26.330 -64.300 -26.160 -63.970 ;
        RECT -32.940 -68.470 -32.770 -64.480 ;
        RECT -32.500 -65.030 -32.330 -64.480 ;
        RECT -26.380 -65.030 -26.210 -64.480 ;
        RECT -26.330 -66.360 -26.160 -66.030 ;
        RECT -32.150 -68.470 -31.980 -66.470 ;
        RECT -26.730 -68.490 -26.560 -66.490 ;
        RECT -32.500 -71.520 -32.330 -68.730 ;
        RECT -26.340 -68.950 -26.170 -68.620 ;
        RECT -25.940 -71.030 -25.770 -64.480 ;
        RECT -32.500 -71.690 -31.980 -71.520 ;
        RECT -32.150 -71.940 -31.980 -71.690 ;
        RECT -25.340 -72.030 -25.170 -64.030 ;
        RECT -24.900 -72.030 -24.730 -64.030 ;
        RECT -24.380 -72.030 -24.210 -63.790 ;
        RECT -23.940 -72.030 -23.770 -64.030 ;
        RECT -23.410 -72.030 -23.240 -64.030 ;
        RECT -22.970 -72.030 -22.800 -63.450 ;
        RECT -12.560 -63.620 -12.390 -63.390 ;
        RECT -12.210 -63.390 -9.450 -63.280 ;
        RECT -2.310 -63.220 -2.140 -59.040 ;
        RECT -1.870 -60.990 -1.700 -59.040 ;
        RECT -1.870 -61.160 -1.660 -60.990 ;
        RECT -1.870 -62.610 -1.700 -61.160 ;
        RECT -1.870 -62.780 -1.660 -62.610 ;
        RECT -1.870 -63.040 -1.700 -62.780 ;
        RECT -0.750 -63.220 -0.580 -59.040 ;
        RECT -0.310 -60.980 -0.140 -59.040 ;
        RECT 0.220 -60.980 0.390 -59.040 ;
        RECT -0.310 -61.150 0.390 -60.980 ;
        RECT -0.310 -62.600 -0.140 -61.150 ;
        RECT 0.220 -62.600 0.390 -61.150 ;
        RECT -0.310 -62.770 -0.120 -62.600 ;
        RECT 0.200 -62.770 0.390 -62.600 ;
        RECT -0.310 -63.040 -0.140 -62.770 ;
        RECT 0.220 -63.040 0.390 -62.770 ;
        RECT -2.310 -63.390 -0.580 -63.220 ;
        RECT 0.660 -63.220 0.830 -59.040 ;
        RECT 1.750 -60.960 1.920 -59.040 ;
        RECT 1.710 -61.130 1.920 -60.960 ;
        RECT 1.750 -62.610 1.920 -61.130 ;
        RECT 1.710 -62.780 1.920 -62.610 ;
        RECT 1.750 -63.040 1.920 -62.780 ;
        RECT 2.190 -63.220 2.360 -59.040 ;
        RECT 2.830 -61.260 3.000 -60.850 ;
        RECT 0.660 -63.280 2.360 -63.220 ;
        RECT -12.210 -63.450 -10.980 -63.390 ;
        RECT -22.220 -63.820 -21.890 -63.650 ;
        RECT -13.470 -63.830 -13.140 -63.660 ;
        RECT -12.560 -63.790 -11.320 -63.620 ;
        RECT -22.450 -72.030 -22.280 -64.030 ;
        RECT -22.010 -72.030 -21.840 -64.030 ;
        RECT -21.050 -64.310 -20.880 -63.980 ;
        RECT -14.510 -64.300 -14.340 -63.970 ;
        RECT -21.440 -68.470 -21.270 -64.480 ;
        RECT -21.000 -65.030 -20.830 -64.480 ;
        RECT -14.560 -65.030 -14.390 -64.480 ;
        RECT -14.510 -66.360 -14.340 -66.030 ;
        RECT -20.650 -68.470 -20.480 -66.470 ;
        RECT -14.910 -68.490 -14.740 -66.490 ;
        RECT -21.000 -71.520 -20.830 -68.730 ;
        RECT -14.520 -68.950 -14.350 -68.620 ;
        RECT -14.120 -71.030 -13.950 -64.480 ;
        RECT -21.000 -71.690 -20.480 -71.520 ;
        RECT -20.650 -71.930 -20.480 -71.690 ;
        RECT -13.520 -72.030 -13.350 -64.030 ;
        RECT -13.080 -72.030 -12.910 -64.030 ;
        RECT -12.560 -72.030 -12.390 -63.790 ;
        RECT -12.120 -72.030 -11.950 -64.030 ;
        RECT -11.590 -72.030 -11.420 -64.030 ;
        RECT -11.150 -72.030 -10.980 -63.450 ;
        RECT -0.750 -63.620 -0.580 -63.390 ;
        RECT -0.400 -63.390 2.360 -63.280 ;
        RECT 9.500 -63.220 9.670 -59.040 ;
        RECT 9.940 -60.990 10.110 -59.040 ;
        RECT 9.940 -61.160 10.150 -60.990 ;
        RECT 9.940 -62.610 10.110 -61.160 ;
        RECT 9.940 -62.780 10.150 -62.610 ;
        RECT 9.940 -63.040 10.110 -62.780 ;
        RECT 11.060 -63.220 11.230 -59.040 ;
        RECT 11.500 -60.980 11.670 -59.040 ;
        RECT 12.030 -60.980 12.200 -59.040 ;
        RECT 11.500 -61.150 12.200 -60.980 ;
        RECT 11.500 -62.600 11.670 -61.150 ;
        RECT 12.030 -62.600 12.200 -61.150 ;
        RECT 11.500 -62.770 11.690 -62.600 ;
        RECT 12.010 -62.770 12.200 -62.600 ;
        RECT 11.500 -63.040 11.670 -62.770 ;
        RECT 12.030 -63.040 12.200 -62.770 ;
        RECT 9.500 -63.390 11.230 -63.220 ;
        RECT 12.470 -63.220 12.640 -59.040 ;
        RECT 13.560 -60.960 13.730 -59.040 ;
        RECT 13.520 -61.130 13.730 -60.960 ;
        RECT 13.560 -62.610 13.730 -61.130 ;
        RECT 13.520 -62.780 13.730 -62.610 ;
        RECT 13.560 -63.040 13.730 -62.780 ;
        RECT 14.000 -63.220 14.170 -59.040 ;
        RECT 14.640 -61.260 14.810 -60.850 ;
        RECT 12.470 -63.280 14.170 -63.220 ;
        RECT -0.400 -63.450 0.830 -63.390 ;
        RECT -10.400 -63.820 -10.070 -63.650 ;
        RECT -1.660 -63.830 -1.330 -63.660 ;
        RECT -0.750 -63.790 0.490 -63.620 ;
        RECT -10.630 -72.030 -10.460 -64.030 ;
        RECT -10.190 -72.030 -10.020 -64.030 ;
        RECT -9.230 -64.310 -9.060 -63.980 ;
        RECT -2.700 -64.300 -2.530 -63.970 ;
        RECT -9.620 -68.470 -9.450 -64.480 ;
        RECT -9.180 -65.030 -9.010 -64.480 ;
        RECT -2.750 -65.030 -2.580 -64.480 ;
        RECT -2.700 -66.360 -2.530 -66.030 ;
        RECT -8.830 -68.470 -8.660 -66.470 ;
        RECT -3.100 -68.490 -2.930 -66.490 ;
        RECT -9.180 -71.520 -9.010 -68.730 ;
        RECT -2.710 -68.950 -2.540 -68.620 ;
        RECT -2.310 -71.030 -2.140 -64.480 ;
        RECT -9.180 -71.690 -8.660 -71.520 ;
        RECT -8.830 -71.930 -8.660 -71.690 ;
        RECT -1.710 -72.030 -1.540 -64.030 ;
        RECT -1.270 -72.030 -1.100 -64.030 ;
        RECT -0.750 -72.030 -0.580 -63.790 ;
        RECT -0.310 -72.030 -0.140 -64.030 ;
        RECT 0.220 -72.030 0.390 -64.030 ;
        RECT 0.660 -72.030 0.830 -63.450 ;
        RECT 11.060 -63.620 11.230 -63.390 ;
        RECT 11.410 -63.390 14.170 -63.280 ;
        RECT 21.320 -63.220 21.490 -59.040 ;
        RECT 21.760 -60.990 21.930 -59.040 ;
        RECT 21.760 -61.160 21.970 -60.990 ;
        RECT 21.760 -62.610 21.930 -61.160 ;
        RECT 21.760 -62.780 21.970 -62.610 ;
        RECT 21.760 -63.040 21.930 -62.780 ;
        RECT 22.880 -63.220 23.050 -59.040 ;
        RECT 23.320 -60.980 23.490 -59.040 ;
        RECT 23.850 -60.980 24.020 -59.040 ;
        RECT 23.320 -61.150 24.020 -60.980 ;
        RECT 23.320 -62.600 23.490 -61.150 ;
        RECT 23.850 -62.600 24.020 -61.150 ;
        RECT 23.320 -62.770 23.510 -62.600 ;
        RECT 23.830 -62.770 24.020 -62.600 ;
        RECT 23.320 -63.040 23.490 -62.770 ;
        RECT 23.850 -63.040 24.020 -62.770 ;
        RECT 21.320 -63.390 23.050 -63.220 ;
        RECT 24.290 -63.220 24.460 -59.040 ;
        RECT 25.380 -60.960 25.550 -59.040 ;
        RECT 25.340 -61.130 25.550 -60.960 ;
        RECT 25.380 -62.610 25.550 -61.130 ;
        RECT 25.340 -62.780 25.550 -62.610 ;
        RECT 25.380 -63.040 25.550 -62.780 ;
        RECT 25.820 -63.220 25.990 -59.040 ;
        RECT 26.460 -61.260 26.630 -60.850 ;
        RECT 24.290 -63.280 25.990 -63.220 ;
        RECT 11.410 -63.450 12.640 -63.390 ;
        RECT 1.410 -63.820 1.740 -63.650 ;
        RECT 10.150 -63.830 10.480 -63.660 ;
        RECT 11.060 -63.790 12.300 -63.620 ;
        RECT 1.180 -72.030 1.350 -64.030 ;
        RECT 1.620 -72.030 1.790 -64.030 ;
        RECT 2.580 -64.310 2.750 -63.980 ;
        RECT 9.110 -64.300 9.280 -63.970 ;
        RECT 2.190 -68.470 2.360 -64.480 ;
        RECT 2.630 -65.030 2.800 -64.480 ;
        RECT 9.060 -65.030 9.230 -64.480 ;
        RECT 9.110 -66.360 9.280 -66.030 ;
        RECT 2.980 -68.470 3.150 -66.470 ;
        RECT 8.710 -68.490 8.880 -66.490 ;
        RECT 2.630 -71.520 2.800 -68.730 ;
        RECT 9.100 -68.950 9.270 -68.620 ;
        RECT 9.500 -71.030 9.670 -64.480 ;
        RECT 2.630 -71.690 3.150 -71.520 ;
        RECT 2.980 -71.930 3.150 -71.690 ;
        RECT 10.100 -72.030 10.270 -64.030 ;
        RECT 10.540 -72.030 10.710 -64.030 ;
        RECT 11.060 -72.030 11.230 -63.790 ;
        RECT 11.500 -72.030 11.670 -64.030 ;
        RECT 12.030 -72.030 12.200 -64.030 ;
        RECT 12.470 -72.030 12.640 -63.450 ;
        RECT 22.880 -63.620 23.050 -63.390 ;
        RECT 23.230 -63.390 25.990 -63.280 ;
        RECT 33.140 -63.220 33.310 -59.040 ;
        RECT 33.580 -60.990 33.750 -59.040 ;
        RECT 33.580 -61.160 33.790 -60.990 ;
        RECT 33.580 -62.610 33.750 -61.160 ;
        RECT 33.580 -62.780 33.790 -62.610 ;
        RECT 33.580 -63.040 33.750 -62.780 ;
        RECT 34.700 -63.220 34.870 -59.040 ;
        RECT 35.140 -60.980 35.310 -59.040 ;
        RECT 35.670 -60.980 35.840 -59.040 ;
        RECT 35.140 -61.150 35.840 -60.980 ;
        RECT 35.140 -62.600 35.310 -61.150 ;
        RECT 35.670 -62.600 35.840 -61.150 ;
        RECT 35.140 -62.770 35.330 -62.600 ;
        RECT 35.650 -62.770 35.840 -62.600 ;
        RECT 35.140 -63.040 35.310 -62.770 ;
        RECT 35.670 -63.040 35.840 -62.770 ;
        RECT 33.140 -63.390 34.870 -63.220 ;
        RECT 36.110 -63.220 36.280 -59.040 ;
        RECT 37.200 -60.960 37.370 -59.040 ;
        RECT 37.160 -61.130 37.370 -60.960 ;
        RECT 37.200 -62.610 37.370 -61.130 ;
        RECT 37.160 -62.780 37.370 -62.610 ;
        RECT 37.200 -63.040 37.370 -62.780 ;
        RECT 37.640 -63.220 37.810 -59.040 ;
        RECT 38.280 -61.260 38.450 -60.850 ;
        RECT 36.110 -63.280 37.810 -63.220 ;
        RECT 23.230 -63.450 24.460 -63.390 ;
        RECT 13.220 -63.820 13.550 -63.650 ;
        RECT 21.970 -63.830 22.300 -63.660 ;
        RECT 22.880 -63.790 24.120 -63.620 ;
        RECT 12.990 -72.030 13.160 -64.030 ;
        RECT 13.430 -72.030 13.600 -64.030 ;
        RECT 14.390 -64.310 14.560 -63.980 ;
        RECT 20.930 -64.300 21.100 -63.970 ;
        RECT 14.000 -68.470 14.170 -64.480 ;
        RECT 14.440 -65.030 14.610 -64.480 ;
        RECT 20.880 -65.030 21.050 -64.480 ;
        RECT 20.930 -66.360 21.100 -66.030 ;
        RECT 14.790 -68.470 14.960 -66.470 ;
        RECT 20.530 -68.490 20.700 -66.490 ;
        RECT 14.440 -71.520 14.610 -68.730 ;
        RECT 20.920 -68.950 21.090 -68.620 ;
        RECT 21.320 -71.030 21.490 -64.480 ;
        RECT 14.440 -71.690 14.960 -71.520 ;
        RECT 14.790 -71.930 14.960 -71.690 ;
        RECT 21.920 -72.030 22.090 -64.030 ;
        RECT 22.360 -72.030 22.530 -64.030 ;
        RECT 22.880 -72.030 23.050 -63.790 ;
        RECT 23.320 -72.030 23.490 -64.030 ;
        RECT 23.850 -72.030 24.020 -64.030 ;
        RECT 24.290 -72.030 24.460 -63.450 ;
        RECT 34.700 -63.620 34.870 -63.390 ;
        RECT 35.050 -63.390 37.810 -63.280 ;
        RECT 44.960 -63.220 45.130 -59.040 ;
        RECT 45.400 -60.990 45.570 -59.040 ;
        RECT 45.400 -61.160 45.610 -60.990 ;
        RECT 45.400 -62.610 45.570 -61.160 ;
        RECT 45.400 -62.780 45.610 -62.610 ;
        RECT 45.400 -63.040 45.570 -62.780 ;
        RECT 46.520 -63.220 46.690 -59.040 ;
        RECT 46.960 -60.980 47.130 -59.040 ;
        RECT 47.490 -60.980 47.660 -59.040 ;
        RECT 46.960 -61.150 47.660 -60.980 ;
        RECT 46.960 -62.600 47.130 -61.150 ;
        RECT 47.490 -62.600 47.660 -61.150 ;
        RECT 46.960 -62.770 47.150 -62.600 ;
        RECT 47.470 -62.770 47.660 -62.600 ;
        RECT 46.960 -63.040 47.130 -62.770 ;
        RECT 47.490 -63.040 47.660 -62.770 ;
        RECT 44.960 -63.390 46.690 -63.220 ;
        RECT 47.930 -63.220 48.100 -59.040 ;
        RECT 49.020 -60.960 49.190 -59.040 ;
        RECT 48.980 -61.130 49.190 -60.960 ;
        RECT 49.020 -62.610 49.190 -61.130 ;
        RECT 48.980 -62.780 49.190 -62.610 ;
        RECT 49.020 -63.040 49.190 -62.780 ;
        RECT 49.460 -63.220 49.630 -59.040 ;
        RECT 50.100 -61.260 50.270 -60.850 ;
        RECT 47.930 -63.280 49.630 -63.220 ;
        RECT 35.050 -63.450 36.280 -63.390 ;
        RECT 25.040 -63.820 25.370 -63.650 ;
        RECT 33.790 -63.830 34.120 -63.660 ;
        RECT 34.700 -63.790 35.940 -63.620 ;
        RECT 24.810 -72.030 24.980 -64.030 ;
        RECT 25.250 -72.030 25.420 -64.030 ;
        RECT 26.210 -64.310 26.380 -63.980 ;
        RECT 32.750 -64.300 32.920 -63.970 ;
        RECT 25.820 -68.470 25.990 -64.480 ;
        RECT 26.260 -65.030 26.430 -64.480 ;
        RECT 32.700 -65.030 32.870 -64.480 ;
        RECT 32.750 -66.360 32.920 -66.030 ;
        RECT 26.610 -68.470 26.780 -66.470 ;
        RECT 32.350 -68.490 32.520 -66.490 ;
        RECT 26.260 -71.520 26.430 -68.730 ;
        RECT 32.740 -68.950 32.910 -68.620 ;
        RECT 33.140 -71.030 33.310 -64.480 ;
        RECT 26.260 -71.690 26.780 -71.520 ;
        RECT 26.610 -71.930 26.780 -71.690 ;
        RECT 33.740 -72.030 33.910 -64.030 ;
        RECT 34.180 -72.030 34.350 -64.030 ;
        RECT 34.700 -72.030 34.870 -63.790 ;
        RECT 35.140 -72.030 35.310 -64.030 ;
        RECT 35.670 -72.030 35.840 -64.030 ;
        RECT 36.110 -72.030 36.280 -63.450 ;
        RECT 46.520 -63.620 46.690 -63.390 ;
        RECT 46.870 -63.390 49.630 -63.280 ;
        RECT 56.780 -63.220 56.950 -59.040 ;
        RECT 57.220 -60.990 57.390 -59.040 ;
        RECT 57.220 -61.160 57.430 -60.990 ;
        RECT 57.220 -62.610 57.390 -61.160 ;
        RECT 57.220 -62.780 57.430 -62.610 ;
        RECT 57.220 -63.040 57.390 -62.780 ;
        RECT 58.340 -63.220 58.510 -59.040 ;
        RECT 58.780 -60.980 58.950 -59.040 ;
        RECT 59.310 -60.980 59.480 -59.040 ;
        RECT 58.780 -61.150 59.480 -60.980 ;
        RECT 58.780 -62.600 58.950 -61.150 ;
        RECT 59.310 -62.600 59.480 -61.150 ;
        RECT 58.780 -62.770 58.970 -62.600 ;
        RECT 59.290 -62.770 59.480 -62.600 ;
        RECT 58.780 -63.040 58.950 -62.770 ;
        RECT 59.310 -63.040 59.480 -62.770 ;
        RECT 56.780 -63.390 58.510 -63.220 ;
        RECT 59.750 -63.220 59.920 -59.040 ;
        RECT 60.840 -60.960 61.010 -59.040 ;
        RECT 60.800 -61.130 61.010 -60.960 ;
        RECT 60.840 -62.610 61.010 -61.130 ;
        RECT 60.800 -62.780 61.010 -62.610 ;
        RECT 60.840 -63.040 61.010 -62.780 ;
        RECT 61.280 -63.220 61.450 -59.040 ;
        RECT 61.920 -61.260 62.090 -60.850 ;
        RECT 59.750 -63.280 61.450 -63.220 ;
        RECT 46.870 -63.450 48.100 -63.390 ;
        RECT 36.860 -63.820 37.190 -63.650 ;
        RECT 45.610 -63.830 45.940 -63.660 ;
        RECT 46.520 -63.790 47.760 -63.620 ;
        RECT 36.630 -72.030 36.800 -64.030 ;
        RECT 37.070 -72.030 37.240 -64.030 ;
        RECT 38.030 -64.310 38.200 -63.980 ;
        RECT 44.570 -64.300 44.740 -63.970 ;
        RECT 37.640 -68.470 37.810 -64.480 ;
        RECT 38.080 -65.030 38.250 -64.480 ;
        RECT 44.520 -65.030 44.690 -64.480 ;
        RECT 44.570 -66.360 44.740 -66.030 ;
        RECT 38.430 -68.470 38.600 -66.470 ;
        RECT 44.170 -68.490 44.340 -66.490 ;
        RECT 38.080 -71.520 38.250 -68.730 ;
        RECT 44.560 -68.950 44.730 -68.620 ;
        RECT 44.960 -71.030 45.130 -64.480 ;
        RECT 38.080 -71.690 38.600 -71.520 ;
        RECT 38.430 -71.930 38.600 -71.690 ;
        RECT 45.560 -72.030 45.730 -64.030 ;
        RECT 46.000 -72.030 46.170 -64.030 ;
        RECT 46.520 -72.030 46.690 -63.790 ;
        RECT 46.960 -72.030 47.130 -64.030 ;
        RECT 47.490 -72.030 47.660 -64.030 ;
        RECT 47.930 -72.030 48.100 -63.450 ;
        RECT 58.340 -63.620 58.510 -63.390 ;
        RECT 58.690 -63.390 61.450 -63.280 ;
        RECT 68.600 -63.220 68.770 -59.040 ;
        RECT 69.040 -60.990 69.210 -59.040 ;
        RECT 69.040 -61.160 69.250 -60.990 ;
        RECT 69.040 -62.610 69.210 -61.160 ;
        RECT 69.040 -62.780 69.250 -62.610 ;
        RECT 69.040 -63.040 69.210 -62.780 ;
        RECT 70.160 -63.220 70.330 -59.040 ;
        RECT 70.600 -60.980 70.770 -59.040 ;
        RECT 71.130 -60.980 71.300 -59.040 ;
        RECT 70.600 -61.150 71.300 -60.980 ;
        RECT 70.600 -62.600 70.770 -61.150 ;
        RECT 71.130 -62.600 71.300 -61.150 ;
        RECT 70.600 -62.770 70.790 -62.600 ;
        RECT 71.110 -62.770 71.300 -62.600 ;
        RECT 70.600 -63.040 70.770 -62.770 ;
        RECT 71.130 -63.040 71.300 -62.770 ;
        RECT 68.600 -63.390 70.330 -63.220 ;
        RECT 71.570 -63.220 71.740 -59.040 ;
        RECT 72.660 -60.960 72.830 -59.040 ;
        RECT 72.620 -61.130 72.830 -60.960 ;
        RECT 72.660 -62.610 72.830 -61.130 ;
        RECT 72.620 -62.780 72.830 -62.610 ;
        RECT 72.660 -63.040 72.830 -62.780 ;
        RECT 73.100 -63.220 73.270 -59.040 ;
        RECT 73.740 -61.260 73.910 -60.850 ;
        RECT 71.570 -63.280 73.270 -63.220 ;
        RECT 58.690 -63.450 59.920 -63.390 ;
        RECT 48.680 -63.820 49.010 -63.650 ;
        RECT 57.430 -63.830 57.760 -63.660 ;
        RECT 58.340 -63.790 59.580 -63.620 ;
        RECT 48.450 -72.030 48.620 -64.030 ;
        RECT 48.890 -72.030 49.060 -64.030 ;
        RECT 49.850 -64.310 50.020 -63.980 ;
        RECT 56.390 -64.300 56.560 -63.970 ;
        RECT 49.460 -68.470 49.630 -64.480 ;
        RECT 49.900 -65.030 50.070 -64.480 ;
        RECT 56.340 -65.030 56.510 -64.480 ;
        RECT 56.390 -66.360 56.560 -66.030 ;
        RECT 50.250 -68.470 50.420 -66.470 ;
        RECT 55.990 -68.490 56.160 -66.490 ;
        RECT 49.900 -71.520 50.070 -68.730 ;
        RECT 56.380 -68.950 56.550 -68.620 ;
        RECT 56.780 -71.030 56.950 -64.480 ;
        RECT 49.900 -71.690 50.420 -71.520 ;
        RECT 50.250 -71.930 50.420 -71.690 ;
        RECT 57.380 -72.030 57.550 -64.030 ;
        RECT 57.820 -72.030 57.990 -64.030 ;
        RECT 58.340 -72.030 58.510 -63.790 ;
        RECT 58.780 -72.030 58.950 -64.030 ;
        RECT 59.310 -72.030 59.480 -64.030 ;
        RECT 59.750 -72.030 59.920 -63.450 ;
        RECT 70.160 -63.620 70.330 -63.390 ;
        RECT 70.510 -63.390 73.270 -63.280 ;
        RECT 80.420 -63.220 80.590 -59.040 ;
        RECT 80.860 -60.990 81.030 -59.040 ;
        RECT 80.860 -61.160 81.070 -60.990 ;
        RECT 80.860 -62.610 81.030 -61.160 ;
        RECT 80.860 -62.780 81.070 -62.610 ;
        RECT 80.860 -63.040 81.030 -62.780 ;
        RECT 81.980 -63.220 82.150 -59.040 ;
        RECT 82.420 -60.980 82.590 -59.040 ;
        RECT 82.950 -60.980 83.120 -59.040 ;
        RECT 82.420 -61.150 83.120 -60.980 ;
        RECT 82.420 -62.600 82.590 -61.150 ;
        RECT 82.950 -62.600 83.120 -61.150 ;
        RECT 82.420 -62.770 82.610 -62.600 ;
        RECT 82.930 -62.770 83.120 -62.600 ;
        RECT 82.420 -63.040 82.590 -62.770 ;
        RECT 82.950 -63.040 83.120 -62.770 ;
        RECT 80.420 -63.390 82.150 -63.220 ;
        RECT 83.390 -63.220 83.560 -59.040 ;
        RECT 84.480 -60.960 84.650 -59.040 ;
        RECT 84.440 -61.130 84.650 -60.960 ;
        RECT 84.480 -62.610 84.650 -61.130 ;
        RECT 84.440 -62.780 84.650 -62.610 ;
        RECT 84.480 -63.040 84.650 -62.780 ;
        RECT 84.920 -63.220 85.090 -59.040 ;
        RECT 85.560 -61.260 85.730 -60.850 ;
        RECT 83.390 -63.280 85.090 -63.220 ;
        RECT 70.510 -63.450 71.740 -63.390 ;
        RECT 60.500 -63.820 60.830 -63.650 ;
        RECT 69.250 -63.830 69.580 -63.660 ;
        RECT 70.160 -63.790 71.400 -63.620 ;
        RECT 60.270 -72.030 60.440 -64.030 ;
        RECT 60.710 -72.030 60.880 -64.030 ;
        RECT 61.670 -64.310 61.840 -63.980 ;
        RECT 68.210 -64.300 68.380 -63.970 ;
        RECT 61.280 -68.470 61.450 -64.480 ;
        RECT 61.720 -65.030 61.890 -64.480 ;
        RECT 68.160 -65.030 68.330 -64.480 ;
        RECT 68.210 -66.360 68.380 -66.030 ;
        RECT 62.070 -68.470 62.240 -66.470 ;
        RECT 67.810 -68.490 67.980 -66.490 ;
        RECT 61.720 -71.520 61.890 -68.730 ;
        RECT 68.200 -68.950 68.370 -68.620 ;
        RECT 68.600 -71.030 68.770 -64.480 ;
        RECT 61.720 -71.690 62.240 -71.520 ;
        RECT 62.070 -71.930 62.240 -71.690 ;
        RECT 69.200 -72.030 69.370 -64.030 ;
        RECT 69.640 -72.030 69.810 -64.030 ;
        RECT 70.160 -72.030 70.330 -63.790 ;
        RECT 70.600 -72.030 70.770 -64.030 ;
        RECT 71.130 -72.030 71.300 -64.030 ;
        RECT 71.570 -72.030 71.740 -63.450 ;
        RECT 81.980 -63.620 82.150 -63.390 ;
        RECT 82.330 -63.390 85.090 -63.280 ;
        RECT 92.260 -63.220 92.430 -59.040 ;
        RECT 92.700 -60.990 92.870 -59.040 ;
        RECT 92.700 -61.160 92.910 -60.990 ;
        RECT 92.700 -62.610 92.870 -61.160 ;
        RECT 92.700 -62.780 92.910 -62.610 ;
        RECT 92.700 -63.040 92.870 -62.780 ;
        RECT 93.820 -63.220 93.990 -59.040 ;
        RECT 94.260 -60.980 94.430 -59.040 ;
        RECT 94.790 -60.980 94.960 -59.040 ;
        RECT 94.260 -61.150 94.960 -60.980 ;
        RECT 94.260 -62.600 94.430 -61.150 ;
        RECT 94.790 -62.600 94.960 -61.150 ;
        RECT 94.260 -62.770 94.450 -62.600 ;
        RECT 94.770 -62.770 94.960 -62.600 ;
        RECT 94.260 -63.040 94.430 -62.770 ;
        RECT 94.790 -63.040 94.960 -62.770 ;
        RECT 92.260 -63.390 93.990 -63.220 ;
        RECT 95.230 -63.220 95.400 -59.040 ;
        RECT 96.320 -60.960 96.490 -59.040 ;
        RECT 96.280 -61.130 96.490 -60.960 ;
        RECT 96.320 -62.610 96.490 -61.130 ;
        RECT 96.280 -62.780 96.490 -62.610 ;
        RECT 96.320 -63.040 96.490 -62.780 ;
        RECT 96.760 -63.220 96.930 -59.040 ;
        RECT 97.400 -61.260 97.570 -60.850 ;
        RECT 95.230 -63.280 96.930 -63.220 ;
        RECT 82.330 -63.450 83.560 -63.390 ;
        RECT 72.320 -63.820 72.650 -63.650 ;
        RECT 81.070 -63.830 81.400 -63.660 ;
        RECT 81.980 -63.790 83.220 -63.620 ;
        RECT 72.090 -72.030 72.260 -64.030 ;
        RECT 72.530 -72.030 72.700 -64.030 ;
        RECT 73.490 -64.310 73.660 -63.980 ;
        RECT 80.030 -64.300 80.200 -63.970 ;
        RECT 73.100 -68.470 73.270 -64.480 ;
        RECT 73.540 -65.030 73.710 -64.480 ;
        RECT 79.980 -65.030 80.150 -64.480 ;
        RECT 80.030 -66.360 80.200 -66.030 ;
        RECT 73.890 -68.470 74.060 -66.470 ;
        RECT 79.630 -68.490 79.800 -66.490 ;
        RECT 73.540 -71.520 73.710 -68.730 ;
        RECT 80.020 -68.950 80.190 -68.620 ;
        RECT 80.420 -71.030 80.590 -64.480 ;
        RECT 73.540 -71.690 74.060 -71.520 ;
        RECT 73.890 -71.930 74.060 -71.690 ;
        RECT 81.020 -72.030 81.190 -64.030 ;
        RECT 81.460 -72.030 81.630 -64.030 ;
        RECT 81.980 -72.030 82.150 -63.790 ;
        RECT 82.420 -72.030 82.590 -64.030 ;
        RECT 82.950 -72.030 83.120 -64.030 ;
        RECT 83.390 -72.030 83.560 -63.450 ;
        RECT 93.820 -63.620 93.990 -63.390 ;
        RECT 94.170 -63.390 96.930 -63.280 ;
        RECT 104.100 -63.220 104.270 -59.040 ;
        RECT 104.540 -60.990 104.710 -59.040 ;
        RECT 104.540 -61.160 104.750 -60.990 ;
        RECT 104.540 -62.610 104.710 -61.160 ;
        RECT 104.540 -62.780 104.750 -62.610 ;
        RECT 104.540 -63.040 104.710 -62.780 ;
        RECT 105.660 -63.220 105.830 -59.040 ;
        RECT 106.100 -60.980 106.270 -59.040 ;
        RECT 106.630 -60.980 106.800 -59.040 ;
        RECT 106.100 -61.150 106.800 -60.980 ;
        RECT 106.100 -62.600 106.270 -61.150 ;
        RECT 106.630 -62.600 106.800 -61.150 ;
        RECT 106.100 -62.770 106.290 -62.600 ;
        RECT 106.610 -62.770 106.800 -62.600 ;
        RECT 106.100 -63.040 106.270 -62.770 ;
        RECT 106.630 -63.040 106.800 -62.770 ;
        RECT 104.100 -63.390 105.830 -63.220 ;
        RECT 107.070 -63.220 107.240 -59.040 ;
        RECT 108.160 -60.960 108.330 -59.040 ;
        RECT 108.120 -61.130 108.330 -60.960 ;
        RECT 108.160 -62.610 108.330 -61.130 ;
        RECT 108.120 -62.780 108.330 -62.610 ;
        RECT 108.160 -63.040 108.330 -62.780 ;
        RECT 108.600 -63.220 108.770 -59.040 ;
        RECT 109.240 -61.260 109.410 -60.850 ;
        RECT 107.070 -63.280 108.770 -63.220 ;
        RECT 94.170 -63.450 95.400 -63.390 ;
        RECT 84.140 -63.820 84.470 -63.650 ;
        RECT 92.910 -63.830 93.240 -63.660 ;
        RECT 93.820 -63.790 95.060 -63.620 ;
        RECT 83.910 -72.030 84.080 -64.030 ;
        RECT 84.350 -72.030 84.520 -64.030 ;
        RECT 85.310 -64.310 85.480 -63.980 ;
        RECT 91.870 -64.300 92.040 -63.970 ;
        RECT 84.920 -68.470 85.090 -64.480 ;
        RECT 85.360 -65.030 85.530 -64.480 ;
        RECT 91.820 -65.030 91.990 -64.480 ;
        RECT 91.870 -66.360 92.040 -66.030 ;
        RECT 85.710 -68.470 85.880 -66.470 ;
        RECT 91.470 -68.490 91.640 -66.490 ;
        RECT 85.360 -71.520 85.530 -68.730 ;
        RECT 91.860 -68.950 92.030 -68.620 ;
        RECT 92.260 -71.030 92.430 -64.480 ;
        RECT 85.360 -71.690 85.880 -71.520 ;
        RECT 85.710 -71.930 85.880 -71.690 ;
        RECT 92.860 -72.030 93.030 -64.030 ;
        RECT 93.300 -72.030 93.470 -64.030 ;
        RECT 93.820 -72.030 93.990 -63.790 ;
        RECT 94.260 -72.030 94.430 -64.030 ;
        RECT 94.790 -72.030 94.960 -64.030 ;
        RECT 95.230 -72.030 95.400 -63.450 ;
        RECT 105.660 -63.620 105.830 -63.390 ;
        RECT 106.010 -63.390 108.770 -63.280 ;
        RECT 115.970 -63.220 116.140 -59.040 ;
        RECT 116.410 -60.990 116.580 -59.040 ;
        RECT 116.410 -61.160 116.620 -60.990 ;
        RECT 116.410 -62.610 116.580 -61.160 ;
        RECT 116.410 -62.780 116.620 -62.610 ;
        RECT 116.410 -63.040 116.580 -62.780 ;
        RECT 117.530 -63.220 117.700 -59.040 ;
        RECT 117.970 -60.980 118.140 -59.040 ;
        RECT 118.500 -60.980 118.670 -59.040 ;
        RECT 117.970 -61.150 118.670 -60.980 ;
        RECT 117.970 -62.600 118.140 -61.150 ;
        RECT 118.500 -62.600 118.670 -61.150 ;
        RECT 117.970 -62.770 118.160 -62.600 ;
        RECT 118.480 -62.770 118.670 -62.600 ;
        RECT 117.970 -63.040 118.140 -62.770 ;
        RECT 118.500 -63.040 118.670 -62.770 ;
        RECT 115.970 -63.390 117.700 -63.220 ;
        RECT 118.940 -63.220 119.110 -59.040 ;
        RECT 120.030 -60.960 120.200 -59.040 ;
        RECT 119.990 -61.130 120.200 -60.960 ;
        RECT 120.030 -62.610 120.200 -61.130 ;
        RECT 119.990 -62.780 120.200 -62.610 ;
        RECT 120.030 -63.040 120.200 -62.780 ;
        RECT 120.470 -63.220 120.640 -59.040 ;
        RECT 121.110 -61.260 121.280 -60.850 ;
        RECT 118.940 -63.280 120.640 -63.220 ;
        RECT 106.010 -63.450 107.240 -63.390 ;
        RECT 95.980 -63.820 96.310 -63.650 ;
        RECT 104.750 -63.830 105.080 -63.660 ;
        RECT 105.660 -63.790 106.900 -63.620 ;
        RECT 95.750 -72.030 95.920 -64.030 ;
        RECT 96.190 -72.030 96.360 -64.030 ;
        RECT 97.150 -64.310 97.320 -63.980 ;
        RECT 103.710 -64.300 103.880 -63.970 ;
        RECT 96.760 -68.470 96.930 -64.480 ;
        RECT 97.200 -65.030 97.370 -64.480 ;
        RECT 103.660 -65.030 103.830 -64.480 ;
        RECT 103.710 -66.360 103.880 -66.030 ;
        RECT 97.550 -68.470 97.720 -66.470 ;
        RECT 103.310 -68.490 103.480 -66.490 ;
        RECT 97.200 -71.520 97.370 -68.730 ;
        RECT 103.700 -68.950 103.870 -68.620 ;
        RECT 104.100 -71.030 104.270 -64.480 ;
        RECT 97.200 -71.690 97.720 -71.520 ;
        RECT 97.550 -71.930 97.720 -71.690 ;
        RECT 104.700 -72.030 104.870 -64.030 ;
        RECT 105.140 -72.030 105.310 -64.030 ;
        RECT 105.660 -72.030 105.830 -63.790 ;
        RECT 106.100 -72.030 106.270 -64.030 ;
        RECT 106.630 -72.030 106.800 -64.030 ;
        RECT 107.070 -72.030 107.240 -63.450 ;
        RECT 117.530 -63.620 117.700 -63.390 ;
        RECT 117.880 -63.390 120.640 -63.280 ;
        RECT 127.840 -63.220 128.010 -59.040 ;
        RECT 128.280 -60.990 128.450 -59.040 ;
        RECT 128.280 -61.160 128.490 -60.990 ;
        RECT 128.280 -62.610 128.450 -61.160 ;
        RECT 128.280 -62.780 128.490 -62.610 ;
        RECT 128.280 -63.040 128.450 -62.780 ;
        RECT 129.400 -63.220 129.570 -59.040 ;
        RECT 129.840 -60.980 130.010 -59.040 ;
        RECT 130.370 -60.980 130.540 -59.040 ;
        RECT 129.840 -61.150 130.540 -60.980 ;
        RECT 129.840 -62.600 130.010 -61.150 ;
        RECT 130.370 -62.600 130.540 -61.150 ;
        RECT 129.840 -62.770 130.030 -62.600 ;
        RECT 130.350 -62.770 130.540 -62.600 ;
        RECT 129.840 -63.040 130.010 -62.770 ;
        RECT 130.370 -63.040 130.540 -62.770 ;
        RECT 127.840 -63.390 129.570 -63.220 ;
        RECT 130.810 -63.220 130.980 -59.040 ;
        RECT 131.900 -60.960 132.070 -59.040 ;
        RECT 131.860 -61.130 132.070 -60.960 ;
        RECT 131.900 -62.610 132.070 -61.130 ;
        RECT 131.860 -62.780 132.070 -62.610 ;
        RECT 131.900 -63.040 132.070 -62.780 ;
        RECT 132.340 -63.220 132.510 -59.040 ;
        RECT 132.980 -61.260 133.150 -60.850 ;
        RECT 130.810 -63.280 132.510 -63.220 ;
        RECT 117.880 -63.450 119.110 -63.390 ;
        RECT 107.820 -63.820 108.150 -63.650 ;
        RECT 116.620 -63.830 116.950 -63.660 ;
        RECT 117.530 -63.790 118.770 -63.620 ;
        RECT 107.590 -72.030 107.760 -64.030 ;
        RECT 108.030 -72.030 108.200 -64.030 ;
        RECT 108.990 -64.310 109.160 -63.980 ;
        RECT 115.580 -64.300 115.750 -63.970 ;
        RECT 108.600 -68.470 108.770 -64.480 ;
        RECT 109.040 -65.030 109.210 -64.480 ;
        RECT 115.530 -65.030 115.700 -64.480 ;
        RECT 115.580 -66.360 115.750 -66.030 ;
        RECT 109.390 -68.470 109.560 -66.470 ;
        RECT 115.180 -68.490 115.350 -66.490 ;
        RECT 109.040 -71.520 109.210 -68.730 ;
        RECT 115.570 -68.950 115.740 -68.620 ;
        RECT 115.970 -71.030 116.140 -64.480 ;
        RECT 109.040 -71.690 109.560 -71.520 ;
        RECT 109.390 -71.930 109.560 -71.690 ;
        RECT 116.570 -72.030 116.740 -64.030 ;
        RECT 117.010 -72.030 117.180 -64.030 ;
        RECT 117.530 -72.030 117.700 -63.790 ;
        RECT 117.970 -72.030 118.140 -64.030 ;
        RECT 118.500 -72.030 118.670 -64.030 ;
        RECT 118.940 -72.030 119.110 -63.450 ;
        RECT 129.400 -63.620 129.570 -63.390 ;
        RECT 129.750 -63.390 132.510 -63.280 ;
        RECT 136.850 -63.220 137.020 -59.040 ;
        RECT 137.290 -60.990 137.460 -59.040 ;
        RECT 137.290 -61.160 137.500 -60.990 ;
        RECT 137.290 -62.610 137.460 -61.160 ;
        RECT 137.290 -62.780 137.500 -62.610 ;
        RECT 137.290 -63.040 137.460 -62.780 ;
        RECT 138.410 -63.220 138.580 -59.040 ;
        RECT 138.850 -60.980 139.020 -59.040 ;
        RECT 139.380 -60.980 139.550 -59.040 ;
        RECT 138.850 -61.150 139.550 -60.980 ;
        RECT 138.850 -62.600 139.020 -61.150 ;
        RECT 139.380 -62.600 139.550 -61.150 ;
        RECT 138.850 -62.770 139.040 -62.600 ;
        RECT 139.360 -62.770 139.550 -62.600 ;
        RECT 138.850 -63.040 139.020 -62.770 ;
        RECT 139.380 -63.040 139.550 -62.770 ;
        RECT 136.850 -63.390 138.580 -63.220 ;
        RECT 139.820 -63.220 139.990 -59.040 ;
        RECT 140.910 -60.960 141.080 -59.040 ;
        RECT 140.870 -61.130 141.080 -60.960 ;
        RECT 140.910 -62.610 141.080 -61.130 ;
        RECT 140.870 -62.780 141.080 -62.610 ;
        RECT 140.910 -63.040 141.080 -62.780 ;
        RECT 141.350 -63.220 141.520 -59.040 ;
        RECT 141.990 -61.260 142.160 -60.850 ;
        RECT 139.820 -63.280 141.520 -63.220 ;
        RECT 129.750 -63.450 130.980 -63.390 ;
        RECT 119.690 -63.820 120.020 -63.650 ;
        RECT 128.490 -63.830 128.820 -63.660 ;
        RECT 129.400 -63.790 130.640 -63.620 ;
        RECT 119.460 -72.030 119.630 -64.030 ;
        RECT 119.900 -72.030 120.070 -64.030 ;
        RECT 120.860 -64.310 121.030 -63.980 ;
        RECT 127.450 -64.300 127.620 -63.970 ;
        RECT 120.470 -68.470 120.640 -64.480 ;
        RECT 120.910 -65.030 121.080 -64.480 ;
        RECT 127.400 -65.030 127.570 -64.480 ;
        RECT 127.450 -66.360 127.620 -66.030 ;
        RECT 121.260 -68.470 121.430 -66.470 ;
        RECT 127.050 -68.490 127.220 -66.490 ;
        RECT 120.910 -71.520 121.080 -68.730 ;
        RECT 127.440 -68.950 127.610 -68.620 ;
        RECT 127.840 -71.030 128.010 -64.480 ;
        RECT 120.910 -71.690 121.430 -71.520 ;
        RECT 121.260 -71.930 121.430 -71.690 ;
        RECT 128.440 -72.030 128.610 -64.030 ;
        RECT 128.880 -72.030 129.050 -64.030 ;
        RECT 129.400 -72.030 129.570 -63.790 ;
        RECT 129.840 -72.030 130.010 -64.030 ;
        RECT 130.370 -72.030 130.540 -64.030 ;
        RECT 130.810 -72.030 130.980 -63.450 ;
        RECT 138.410 -63.620 138.580 -63.390 ;
        RECT 138.760 -63.390 141.520 -63.280 ;
        RECT 138.760 -63.450 139.990 -63.390 ;
        RECT 131.560 -63.820 131.890 -63.650 ;
        RECT 137.500 -63.830 137.830 -63.660 ;
        RECT 138.410 -63.790 139.650 -63.620 ;
        RECT 131.330 -72.030 131.500 -64.030 ;
        RECT 131.770 -72.030 131.940 -64.030 ;
        RECT 132.730 -64.310 132.900 -63.980 ;
        RECT 136.460 -64.300 136.630 -63.970 ;
        RECT 132.340 -68.470 132.510 -64.480 ;
        RECT 132.780 -65.030 132.950 -64.480 ;
        RECT 136.410 -65.030 136.580 -64.480 ;
        RECT 136.460 -66.360 136.630 -66.030 ;
        RECT 133.130 -68.470 133.300 -66.470 ;
        RECT 136.060 -68.490 136.230 -66.490 ;
        RECT 132.780 -71.520 132.950 -68.730 ;
        RECT 136.450 -68.950 136.620 -68.620 ;
        RECT 136.850 -71.030 137.020 -64.480 ;
        RECT 132.780 -71.690 133.300 -71.520 ;
        RECT 133.130 -71.930 133.300 -71.690 ;
        RECT 137.450 -72.030 137.620 -64.030 ;
        RECT 137.890 -72.030 138.060 -64.030 ;
        RECT 138.410 -72.030 138.580 -63.790 ;
        RECT 138.850 -72.030 139.020 -64.030 ;
        RECT 139.380 -72.030 139.550 -64.030 ;
        RECT 139.820 -72.030 139.990 -63.450 ;
        RECT 140.570 -63.820 140.900 -63.650 ;
        RECT 140.340 -72.030 140.510 -64.030 ;
        RECT 140.780 -72.030 140.950 -64.030 ;
        RECT 141.740 -64.310 141.910 -63.980 ;
        RECT 141.350 -68.470 141.520 -64.480 ;
        RECT 141.790 -65.030 141.960 -64.480 ;
        RECT 142.140 -68.470 142.310 -66.470 ;
        RECT 141.790 -71.520 141.960 -68.730 ;
        RECT 141.790 -71.690 142.310 -71.520 ;
        RECT 142.140 -71.930 142.310 -71.690 ;
        RECT -32.870 -72.630 -32.700 -72.220 ;
        RECT -21.370 -72.630 -21.200 -72.220 ;
        RECT -9.550 -72.630 -9.380 -72.220 ;
        RECT 2.260 -72.630 2.430 -72.220 ;
        RECT 14.070 -72.630 14.240 -72.220 ;
        RECT 25.890 -72.630 26.060 -72.220 ;
        RECT 37.710 -72.630 37.880 -72.220 ;
        RECT 49.530 -72.630 49.700 -72.220 ;
        RECT 61.350 -72.630 61.520 -72.220 ;
        RECT 73.170 -72.630 73.340 -72.220 ;
        RECT 84.990 -72.630 85.160 -72.220 ;
        RECT 96.830 -72.630 97.000 -72.220 ;
        RECT 108.670 -72.630 108.840 -72.220 ;
        RECT 120.540 -72.630 120.710 -72.220 ;
        RECT 132.410 -72.630 132.580 -72.220 ;
        RECT 141.420 -72.630 141.590 -72.220 ;
        RECT -37.840 -76.120 -37.670 -75.790 ;
        RECT -38.230 -78.250 -38.060 -76.250 ;
        RECT -37.880 -80.260 -37.710 -79.710 ;
        RECT -37.440 -80.260 -37.270 -73.710 ;
        RECT -37.830 -80.770 -37.660 -80.440 ;
        RECT -36.840 -80.710 -36.670 -72.710 ;
        RECT -36.400 -80.710 -36.230 -72.710 ;
        RECT -36.790 -81.080 -36.460 -80.910 ;
        RECT -35.880 -80.950 -35.710 -72.710 ;
        RECT -35.440 -80.710 -35.270 -72.710 ;
        RECT -34.910 -80.710 -34.740 -72.710 ;
        RECT -35.880 -81.120 -34.640 -80.950 ;
        RECT -35.880 -81.350 -35.710 -81.120 ;
        RECT -34.470 -81.290 -34.300 -72.710 ;
        RECT -33.950 -80.710 -33.780 -72.710 ;
        RECT -33.510 -80.710 -33.340 -72.710 ;
        RECT -32.150 -73.040 -31.980 -72.740 ;
        RECT -32.500 -73.210 -31.980 -73.040 ;
        RECT -32.500 -76.150 -32.330 -73.210 ;
        RECT -26.340 -76.120 -26.170 -75.790 ;
        RECT -32.940 -80.260 -32.770 -76.270 ;
        RECT -32.150 -78.270 -31.980 -76.270 ;
        RECT -26.730 -78.250 -26.560 -76.250 ;
        RECT -32.500 -80.260 -32.330 -79.710 ;
        RECT -26.380 -80.260 -26.210 -79.710 ;
        RECT -25.940 -80.260 -25.770 -73.710 ;
        RECT -32.550 -80.760 -32.380 -80.430 ;
        RECT -26.330 -80.770 -26.160 -80.440 ;
        RECT -25.340 -80.710 -25.170 -72.710 ;
        RECT -24.900 -80.710 -24.730 -72.710 ;
        RECT -33.720 -81.090 -33.390 -80.920 ;
        RECT -25.290 -81.080 -24.960 -80.910 ;
        RECT -24.380 -80.950 -24.210 -72.710 ;
        RECT -23.940 -80.710 -23.770 -72.710 ;
        RECT -23.410 -80.710 -23.240 -72.710 ;
        RECT -37.440 -81.520 -35.710 -81.350 ;
        RECT -35.530 -81.350 -34.300 -81.290 ;
        RECT -24.380 -81.120 -23.140 -80.950 ;
        RECT -24.380 -81.350 -24.210 -81.120 ;
        RECT -22.970 -81.290 -22.800 -72.710 ;
        RECT -22.450 -80.710 -22.280 -72.710 ;
        RECT -22.010 -80.710 -21.840 -72.710 ;
        RECT -20.650 -73.040 -20.480 -72.730 ;
        RECT -21.000 -73.210 -20.480 -73.040 ;
        RECT -21.000 -76.150 -20.830 -73.210 ;
        RECT -14.520 -76.120 -14.350 -75.790 ;
        RECT -21.440 -80.260 -21.270 -76.270 ;
        RECT -20.650 -78.270 -20.480 -76.270 ;
        RECT -14.910 -78.250 -14.740 -76.250 ;
        RECT -21.000 -80.260 -20.830 -79.710 ;
        RECT -14.560 -80.260 -14.390 -79.710 ;
        RECT -14.120 -80.260 -13.950 -73.710 ;
        RECT -21.050 -80.760 -20.880 -80.430 ;
        RECT -14.510 -80.770 -14.340 -80.440 ;
        RECT -13.520 -80.710 -13.350 -72.710 ;
        RECT -13.080 -80.710 -12.910 -72.710 ;
        RECT -22.220 -81.090 -21.890 -80.920 ;
        RECT -13.470 -81.080 -13.140 -80.910 ;
        RECT -12.560 -80.950 -12.390 -72.710 ;
        RECT -12.120 -80.710 -11.950 -72.710 ;
        RECT -11.590 -80.710 -11.420 -72.710 ;
        RECT -35.530 -81.460 -32.770 -81.350 ;
        RECT -37.440 -85.700 -37.270 -81.520 ;
        RECT -37.000 -81.960 -36.830 -81.700 ;
        RECT -37.000 -82.130 -36.790 -81.960 ;
        RECT -37.000 -83.580 -36.830 -82.130 ;
        RECT -37.000 -83.750 -36.790 -83.580 ;
        RECT -37.000 -85.700 -36.830 -83.750 ;
        RECT -35.880 -85.700 -35.710 -81.520 ;
        RECT -34.470 -81.520 -32.770 -81.460 ;
        RECT -35.440 -81.970 -35.270 -81.700 ;
        RECT -34.910 -81.970 -34.740 -81.700 ;
        RECT -35.440 -82.140 -35.250 -81.970 ;
        RECT -34.930 -82.140 -34.740 -81.970 ;
        RECT -35.440 -83.590 -35.270 -82.140 ;
        RECT -34.910 -83.590 -34.740 -82.140 ;
        RECT -35.440 -83.760 -34.740 -83.590 ;
        RECT -35.440 -85.700 -35.270 -83.760 ;
        RECT -34.910 -85.700 -34.740 -83.760 ;
        RECT -34.470 -85.700 -34.300 -81.520 ;
        RECT -33.380 -81.960 -33.210 -81.700 ;
        RECT -33.420 -82.130 -33.210 -81.960 ;
        RECT -33.380 -83.610 -33.210 -82.130 ;
        RECT -33.420 -83.780 -33.210 -83.610 ;
        RECT -33.380 -85.700 -33.210 -83.780 ;
        RECT -32.940 -85.700 -32.770 -81.520 ;
        RECT -25.940 -81.520 -24.210 -81.350 ;
        RECT -24.030 -81.350 -22.800 -81.290 ;
        RECT -12.560 -81.120 -11.320 -80.950 ;
        RECT -12.560 -81.350 -12.390 -81.120 ;
        RECT -11.150 -81.290 -10.980 -72.710 ;
        RECT -10.630 -80.710 -10.460 -72.710 ;
        RECT -10.190 -80.710 -10.020 -72.710 ;
        RECT -8.830 -73.040 -8.660 -72.730 ;
        RECT -9.180 -73.210 -8.660 -73.040 ;
        RECT -9.180 -76.150 -9.010 -73.210 ;
        RECT -2.710 -76.120 -2.540 -75.790 ;
        RECT -9.620 -80.260 -9.450 -76.270 ;
        RECT -8.830 -78.270 -8.660 -76.270 ;
        RECT -3.100 -78.250 -2.930 -76.250 ;
        RECT -9.180 -80.260 -9.010 -79.710 ;
        RECT -2.750 -80.260 -2.580 -79.710 ;
        RECT -2.310 -80.260 -2.140 -73.710 ;
        RECT -9.230 -80.760 -9.060 -80.430 ;
        RECT -2.700 -80.770 -2.530 -80.440 ;
        RECT -1.710 -80.710 -1.540 -72.710 ;
        RECT -1.270 -80.710 -1.100 -72.710 ;
        RECT -10.400 -81.090 -10.070 -80.920 ;
        RECT -1.660 -81.080 -1.330 -80.910 ;
        RECT -0.750 -80.950 -0.580 -72.710 ;
        RECT -0.310 -80.710 -0.140 -72.710 ;
        RECT 0.220 -80.710 0.390 -72.710 ;
        RECT -24.030 -81.460 -21.270 -81.350 ;
        RECT -32.340 -83.880 -32.170 -83.470 ;
        RECT -25.940 -85.700 -25.770 -81.520 ;
        RECT -25.500 -81.960 -25.330 -81.700 ;
        RECT -25.500 -82.130 -25.290 -81.960 ;
        RECT -25.500 -83.580 -25.330 -82.130 ;
        RECT -25.500 -83.750 -25.290 -83.580 ;
        RECT -25.500 -85.700 -25.330 -83.750 ;
        RECT -24.380 -85.700 -24.210 -81.520 ;
        RECT -22.970 -81.520 -21.270 -81.460 ;
        RECT -23.940 -81.970 -23.770 -81.700 ;
        RECT -23.410 -81.970 -23.240 -81.700 ;
        RECT -23.940 -82.140 -23.750 -81.970 ;
        RECT -23.430 -82.140 -23.240 -81.970 ;
        RECT -23.940 -83.590 -23.770 -82.140 ;
        RECT -23.410 -83.590 -23.240 -82.140 ;
        RECT -23.940 -83.760 -23.240 -83.590 ;
        RECT -23.940 -85.700 -23.770 -83.760 ;
        RECT -23.410 -85.700 -23.240 -83.760 ;
        RECT -22.970 -85.700 -22.800 -81.520 ;
        RECT -21.880 -81.960 -21.710 -81.700 ;
        RECT -21.920 -82.130 -21.710 -81.960 ;
        RECT -21.880 -83.610 -21.710 -82.130 ;
        RECT -21.920 -83.780 -21.710 -83.610 ;
        RECT -21.880 -85.700 -21.710 -83.780 ;
        RECT -21.440 -85.700 -21.270 -81.520 ;
        RECT -14.120 -81.520 -12.390 -81.350 ;
        RECT -12.210 -81.350 -10.980 -81.290 ;
        RECT -0.750 -81.120 0.490 -80.950 ;
        RECT -0.750 -81.350 -0.580 -81.120 ;
        RECT 0.660 -81.290 0.830 -72.710 ;
        RECT 1.180 -80.710 1.350 -72.710 ;
        RECT 1.620 -80.710 1.790 -72.710 ;
        RECT 2.980 -73.040 3.150 -72.730 ;
        RECT 2.630 -73.210 3.150 -73.040 ;
        RECT 2.630 -76.150 2.800 -73.210 ;
        RECT 9.100 -76.120 9.270 -75.790 ;
        RECT 2.190 -80.260 2.360 -76.270 ;
        RECT 2.980 -78.270 3.150 -76.270 ;
        RECT 8.710 -78.250 8.880 -76.250 ;
        RECT 2.630 -80.260 2.800 -79.710 ;
        RECT 9.060 -80.260 9.230 -79.710 ;
        RECT 9.500 -80.260 9.670 -73.710 ;
        RECT 2.580 -80.760 2.750 -80.430 ;
        RECT 9.110 -80.770 9.280 -80.440 ;
        RECT 10.100 -80.710 10.270 -72.710 ;
        RECT 10.540 -80.710 10.710 -72.710 ;
        RECT 1.410 -81.090 1.740 -80.920 ;
        RECT 10.150 -81.080 10.480 -80.910 ;
        RECT 11.060 -80.950 11.230 -72.710 ;
        RECT 11.500 -80.710 11.670 -72.710 ;
        RECT 12.030 -80.710 12.200 -72.710 ;
        RECT -12.210 -81.460 -9.450 -81.350 ;
        RECT -20.840 -83.880 -20.670 -83.470 ;
        RECT -14.120 -85.700 -13.950 -81.520 ;
        RECT -13.680 -81.960 -13.510 -81.700 ;
        RECT -13.680 -82.130 -13.470 -81.960 ;
        RECT -13.680 -83.580 -13.510 -82.130 ;
        RECT -13.680 -83.750 -13.470 -83.580 ;
        RECT -13.680 -85.700 -13.510 -83.750 ;
        RECT -12.560 -85.700 -12.390 -81.520 ;
        RECT -11.150 -81.520 -9.450 -81.460 ;
        RECT -12.120 -81.970 -11.950 -81.700 ;
        RECT -11.590 -81.970 -11.420 -81.700 ;
        RECT -12.120 -82.140 -11.930 -81.970 ;
        RECT -11.610 -82.140 -11.420 -81.970 ;
        RECT -12.120 -83.590 -11.950 -82.140 ;
        RECT -11.590 -83.590 -11.420 -82.140 ;
        RECT -12.120 -83.760 -11.420 -83.590 ;
        RECT -12.120 -85.700 -11.950 -83.760 ;
        RECT -11.590 -85.700 -11.420 -83.760 ;
        RECT -11.150 -85.700 -10.980 -81.520 ;
        RECT -10.060 -81.960 -9.890 -81.700 ;
        RECT -10.100 -82.130 -9.890 -81.960 ;
        RECT -10.060 -83.610 -9.890 -82.130 ;
        RECT -10.100 -83.780 -9.890 -83.610 ;
        RECT -10.060 -85.700 -9.890 -83.780 ;
        RECT -9.620 -85.700 -9.450 -81.520 ;
        RECT -2.310 -81.520 -0.580 -81.350 ;
        RECT -0.400 -81.350 0.830 -81.290 ;
        RECT 11.060 -81.120 12.300 -80.950 ;
        RECT 11.060 -81.350 11.230 -81.120 ;
        RECT 12.470 -81.290 12.640 -72.710 ;
        RECT 12.990 -80.710 13.160 -72.710 ;
        RECT 13.430 -80.710 13.600 -72.710 ;
        RECT 14.790 -73.040 14.960 -72.730 ;
        RECT 14.440 -73.210 14.960 -73.040 ;
        RECT 14.440 -76.150 14.610 -73.210 ;
        RECT 20.920 -76.120 21.090 -75.790 ;
        RECT 14.000 -80.260 14.170 -76.270 ;
        RECT 14.790 -78.270 14.960 -76.270 ;
        RECT 20.530 -78.250 20.700 -76.250 ;
        RECT 14.440 -80.260 14.610 -79.710 ;
        RECT 20.880 -80.260 21.050 -79.710 ;
        RECT 21.320 -80.260 21.490 -73.710 ;
        RECT 14.390 -80.760 14.560 -80.430 ;
        RECT 20.930 -80.770 21.100 -80.440 ;
        RECT 21.920 -80.710 22.090 -72.710 ;
        RECT 22.360 -80.710 22.530 -72.710 ;
        RECT 13.220 -81.090 13.550 -80.920 ;
        RECT 21.970 -81.080 22.300 -80.910 ;
        RECT 22.880 -80.950 23.050 -72.710 ;
        RECT 23.320 -80.710 23.490 -72.710 ;
        RECT 23.850 -80.710 24.020 -72.710 ;
        RECT -0.400 -81.460 2.360 -81.350 ;
        RECT -9.020 -83.880 -8.850 -83.470 ;
        RECT -2.310 -85.700 -2.140 -81.520 ;
        RECT -1.870 -81.960 -1.700 -81.700 ;
        RECT -1.870 -82.130 -1.660 -81.960 ;
        RECT -1.870 -83.580 -1.700 -82.130 ;
        RECT -1.870 -83.750 -1.660 -83.580 ;
        RECT -1.870 -85.700 -1.700 -83.750 ;
        RECT -0.750 -85.700 -0.580 -81.520 ;
        RECT 0.660 -81.520 2.360 -81.460 ;
        RECT -0.310 -81.970 -0.140 -81.700 ;
        RECT 0.220 -81.970 0.390 -81.700 ;
        RECT -0.310 -82.140 -0.120 -81.970 ;
        RECT 0.200 -82.140 0.390 -81.970 ;
        RECT -0.310 -83.590 -0.140 -82.140 ;
        RECT 0.220 -83.590 0.390 -82.140 ;
        RECT -0.310 -83.760 0.390 -83.590 ;
        RECT -0.310 -85.700 -0.140 -83.760 ;
        RECT 0.220 -85.700 0.390 -83.760 ;
        RECT 0.660 -85.700 0.830 -81.520 ;
        RECT 1.750 -81.960 1.920 -81.700 ;
        RECT 1.710 -82.130 1.920 -81.960 ;
        RECT 1.750 -83.610 1.920 -82.130 ;
        RECT 1.710 -83.780 1.920 -83.610 ;
        RECT 1.750 -85.700 1.920 -83.780 ;
        RECT 2.190 -85.700 2.360 -81.520 ;
        RECT 9.500 -81.520 11.230 -81.350 ;
        RECT 11.410 -81.350 12.640 -81.290 ;
        RECT 22.880 -81.120 24.120 -80.950 ;
        RECT 22.880 -81.350 23.050 -81.120 ;
        RECT 24.290 -81.290 24.460 -72.710 ;
        RECT 24.810 -80.710 24.980 -72.710 ;
        RECT 25.250 -80.710 25.420 -72.710 ;
        RECT 26.610 -73.040 26.780 -72.730 ;
        RECT 26.260 -73.210 26.780 -73.040 ;
        RECT 26.260 -76.150 26.430 -73.210 ;
        RECT 32.740 -76.120 32.910 -75.790 ;
        RECT 25.820 -80.260 25.990 -76.270 ;
        RECT 26.610 -78.270 26.780 -76.270 ;
        RECT 32.350 -78.250 32.520 -76.250 ;
        RECT 26.260 -80.260 26.430 -79.710 ;
        RECT 32.700 -80.260 32.870 -79.710 ;
        RECT 33.140 -80.260 33.310 -73.710 ;
        RECT 26.210 -80.760 26.380 -80.430 ;
        RECT 32.750 -80.770 32.920 -80.440 ;
        RECT 33.740 -80.710 33.910 -72.710 ;
        RECT 34.180 -80.710 34.350 -72.710 ;
        RECT 25.040 -81.090 25.370 -80.920 ;
        RECT 33.790 -81.080 34.120 -80.910 ;
        RECT 34.700 -80.950 34.870 -72.710 ;
        RECT 35.140 -80.710 35.310 -72.710 ;
        RECT 35.670 -80.710 35.840 -72.710 ;
        RECT 11.410 -81.460 14.170 -81.350 ;
        RECT 2.790 -83.880 2.960 -83.470 ;
        RECT 9.500 -85.700 9.670 -81.520 ;
        RECT 9.940 -81.960 10.110 -81.700 ;
        RECT 9.940 -82.130 10.150 -81.960 ;
        RECT 9.940 -83.580 10.110 -82.130 ;
        RECT 9.940 -83.750 10.150 -83.580 ;
        RECT 9.940 -85.700 10.110 -83.750 ;
        RECT 11.060 -85.700 11.230 -81.520 ;
        RECT 12.470 -81.520 14.170 -81.460 ;
        RECT 11.500 -81.970 11.670 -81.700 ;
        RECT 12.030 -81.970 12.200 -81.700 ;
        RECT 11.500 -82.140 11.690 -81.970 ;
        RECT 12.010 -82.140 12.200 -81.970 ;
        RECT 11.500 -83.590 11.670 -82.140 ;
        RECT 12.030 -83.590 12.200 -82.140 ;
        RECT 11.500 -83.760 12.200 -83.590 ;
        RECT 11.500 -85.700 11.670 -83.760 ;
        RECT 12.030 -85.700 12.200 -83.760 ;
        RECT 12.470 -85.700 12.640 -81.520 ;
        RECT 13.560 -81.960 13.730 -81.700 ;
        RECT 13.520 -82.130 13.730 -81.960 ;
        RECT 13.560 -83.610 13.730 -82.130 ;
        RECT 13.520 -83.780 13.730 -83.610 ;
        RECT 13.560 -85.700 13.730 -83.780 ;
        RECT 14.000 -85.700 14.170 -81.520 ;
        RECT 21.320 -81.520 23.050 -81.350 ;
        RECT 23.230 -81.350 24.460 -81.290 ;
        RECT 34.700 -81.120 35.940 -80.950 ;
        RECT 34.700 -81.350 34.870 -81.120 ;
        RECT 36.110 -81.290 36.280 -72.710 ;
        RECT 36.630 -80.710 36.800 -72.710 ;
        RECT 37.070 -80.710 37.240 -72.710 ;
        RECT 38.430 -73.040 38.600 -72.730 ;
        RECT 38.080 -73.210 38.600 -73.040 ;
        RECT 38.080 -76.150 38.250 -73.210 ;
        RECT 44.560 -76.120 44.730 -75.790 ;
        RECT 37.640 -80.260 37.810 -76.270 ;
        RECT 38.430 -78.270 38.600 -76.270 ;
        RECT 44.170 -78.250 44.340 -76.250 ;
        RECT 38.080 -80.260 38.250 -79.710 ;
        RECT 44.520 -80.260 44.690 -79.710 ;
        RECT 44.960 -80.260 45.130 -73.710 ;
        RECT 38.030 -80.760 38.200 -80.430 ;
        RECT 44.570 -80.770 44.740 -80.440 ;
        RECT 45.560 -80.710 45.730 -72.710 ;
        RECT 46.000 -80.710 46.170 -72.710 ;
        RECT 36.860 -81.090 37.190 -80.920 ;
        RECT 45.610 -81.080 45.940 -80.910 ;
        RECT 46.520 -80.950 46.690 -72.710 ;
        RECT 46.960 -80.710 47.130 -72.710 ;
        RECT 47.490 -80.710 47.660 -72.710 ;
        RECT 23.230 -81.460 25.990 -81.350 ;
        RECT 14.600 -83.880 14.770 -83.470 ;
        RECT 21.320 -85.700 21.490 -81.520 ;
        RECT 21.760 -81.960 21.930 -81.700 ;
        RECT 21.760 -82.130 21.970 -81.960 ;
        RECT 21.760 -83.580 21.930 -82.130 ;
        RECT 21.760 -83.750 21.970 -83.580 ;
        RECT 21.760 -85.700 21.930 -83.750 ;
        RECT 22.880 -85.700 23.050 -81.520 ;
        RECT 24.290 -81.520 25.990 -81.460 ;
        RECT 23.320 -81.970 23.490 -81.700 ;
        RECT 23.850 -81.970 24.020 -81.700 ;
        RECT 23.320 -82.140 23.510 -81.970 ;
        RECT 23.830 -82.140 24.020 -81.970 ;
        RECT 23.320 -83.590 23.490 -82.140 ;
        RECT 23.850 -83.590 24.020 -82.140 ;
        RECT 23.320 -83.760 24.020 -83.590 ;
        RECT 23.320 -85.700 23.490 -83.760 ;
        RECT 23.850 -85.700 24.020 -83.760 ;
        RECT 24.290 -85.700 24.460 -81.520 ;
        RECT 25.380 -81.960 25.550 -81.700 ;
        RECT 25.340 -82.130 25.550 -81.960 ;
        RECT 25.380 -83.610 25.550 -82.130 ;
        RECT 25.340 -83.780 25.550 -83.610 ;
        RECT 25.380 -85.700 25.550 -83.780 ;
        RECT 25.820 -85.700 25.990 -81.520 ;
        RECT 33.140 -81.520 34.870 -81.350 ;
        RECT 35.050 -81.350 36.280 -81.290 ;
        RECT 46.520 -81.120 47.760 -80.950 ;
        RECT 46.520 -81.350 46.690 -81.120 ;
        RECT 47.930 -81.290 48.100 -72.710 ;
        RECT 48.450 -80.710 48.620 -72.710 ;
        RECT 48.890 -80.710 49.060 -72.710 ;
        RECT 50.250 -73.040 50.420 -72.730 ;
        RECT 49.900 -73.210 50.420 -73.040 ;
        RECT 49.900 -76.150 50.070 -73.210 ;
        RECT 56.380 -76.120 56.550 -75.790 ;
        RECT 49.460 -80.260 49.630 -76.270 ;
        RECT 50.250 -78.270 50.420 -76.270 ;
        RECT 55.990 -78.250 56.160 -76.250 ;
        RECT 49.900 -80.260 50.070 -79.710 ;
        RECT 56.340 -80.260 56.510 -79.710 ;
        RECT 56.780 -80.260 56.950 -73.710 ;
        RECT 49.850 -80.760 50.020 -80.430 ;
        RECT 56.390 -80.770 56.560 -80.440 ;
        RECT 57.380 -80.710 57.550 -72.710 ;
        RECT 57.820 -80.710 57.990 -72.710 ;
        RECT 48.680 -81.090 49.010 -80.920 ;
        RECT 57.430 -81.080 57.760 -80.910 ;
        RECT 58.340 -80.950 58.510 -72.710 ;
        RECT 58.780 -80.710 58.950 -72.710 ;
        RECT 59.310 -80.710 59.480 -72.710 ;
        RECT 35.050 -81.460 37.810 -81.350 ;
        RECT 26.420 -83.880 26.590 -83.470 ;
        RECT 33.140 -85.700 33.310 -81.520 ;
        RECT 33.580 -81.960 33.750 -81.700 ;
        RECT 33.580 -82.130 33.790 -81.960 ;
        RECT 33.580 -83.580 33.750 -82.130 ;
        RECT 33.580 -83.750 33.790 -83.580 ;
        RECT 33.580 -85.700 33.750 -83.750 ;
        RECT 34.700 -85.700 34.870 -81.520 ;
        RECT 36.110 -81.520 37.810 -81.460 ;
        RECT 35.140 -81.970 35.310 -81.700 ;
        RECT 35.670 -81.970 35.840 -81.700 ;
        RECT 35.140 -82.140 35.330 -81.970 ;
        RECT 35.650 -82.140 35.840 -81.970 ;
        RECT 35.140 -83.590 35.310 -82.140 ;
        RECT 35.670 -83.590 35.840 -82.140 ;
        RECT 35.140 -83.760 35.840 -83.590 ;
        RECT 35.140 -85.700 35.310 -83.760 ;
        RECT 35.670 -85.700 35.840 -83.760 ;
        RECT 36.110 -85.700 36.280 -81.520 ;
        RECT 37.200 -81.960 37.370 -81.700 ;
        RECT 37.160 -82.130 37.370 -81.960 ;
        RECT 37.200 -83.610 37.370 -82.130 ;
        RECT 37.160 -83.780 37.370 -83.610 ;
        RECT 37.200 -85.700 37.370 -83.780 ;
        RECT 37.640 -85.700 37.810 -81.520 ;
        RECT 44.960 -81.520 46.690 -81.350 ;
        RECT 46.870 -81.350 48.100 -81.290 ;
        RECT 58.340 -81.120 59.580 -80.950 ;
        RECT 58.340 -81.350 58.510 -81.120 ;
        RECT 59.750 -81.290 59.920 -72.710 ;
        RECT 60.270 -80.710 60.440 -72.710 ;
        RECT 60.710 -80.710 60.880 -72.710 ;
        RECT 62.070 -73.040 62.240 -72.730 ;
        RECT 61.720 -73.210 62.240 -73.040 ;
        RECT 61.720 -76.150 61.890 -73.210 ;
        RECT 68.200 -76.120 68.370 -75.790 ;
        RECT 61.280 -80.260 61.450 -76.270 ;
        RECT 62.070 -78.270 62.240 -76.270 ;
        RECT 67.810 -78.250 67.980 -76.250 ;
        RECT 61.720 -80.260 61.890 -79.710 ;
        RECT 68.160 -80.260 68.330 -79.710 ;
        RECT 68.600 -80.260 68.770 -73.710 ;
        RECT 61.670 -80.760 61.840 -80.430 ;
        RECT 68.210 -80.770 68.380 -80.440 ;
        RECT 69.200 -80.710 69.370 -72.710 ;
        RECT 69.640 -80.710 69.810 -72.710 ;
        RECT 60.500 -81.090 60.830 -80.920 ;
        RECT 69.250 -81.080 69.580 -80.910 ;
        RECT 70.160 -80.950 70.330 -72.710 ;
        RECT 70.600 -80.710 70.770 -72.710 ;
        RECT 71.130 -80.710 71.300 -72.710 ;
        RECT 46.870 -81.460 49.630 -81.350 ;
        RECT 38.240 -83.880 38.410 -83.470 ;
        RECT 44.960 -85.700 45.130 -81.520 ;
        RECT 45.400 -81.960 45.570 -81.700 ;
        RECT 45.400 -82.130 45.610 -81.960 ;
        RECT 45.400 -83.580 45.570 -82.130 ;
        RECT 45.400 -83.750 45.610 -83.580 ;
        RECT 45.400 -85.700 45.570 -83.750 ;
        RECT 46.520 -85.700 46.690 -81.520 ;
        RECT 47.930 -81.520 49.630 -81.460 ;
        RECT 46.960 -81.970 47.130 -81.700 ;
        RECT 47.490 -81.970 47.660 -81.700 ;
        RECT 46.960 -82.140 47.150 -81.970 ;
        RECT 47.470 -82.140 47.660 -81.970 ;
        RECT 46.960 -83.590 47.130 -82.140 ;
        RECT 47.490 -83.590 47.660 -82.140 ;
        RECT 46.960 -83.760 47.660 -83.590 ;
        RECT 46.960 -85.700 47.130 -83.760 ;
        RECT 47.490 -85.700 47.660 -83.760 ;
        RECT 47.930 -85.700 48.100 -81.520 ;
        RECT 49.020 -81.960 49.190 -81.700 ;
        RECT 48.980 -82.130 49.190 -81.960 ;
        RECT 49.020 -83.610 49.190 -82.130 ;
        RECT 48.980 -83.780 49.190 -83.610 ;
        RECT 49.020 -85.700 49.190 -83.780 ;
        RECT 49.460 -85.700 49.630 -81.520 ;
        RECT 56.780 -81.520 58.510 -81.350 ;
        RECT 58.690 -81.350 59.920 -81.290 ;
        RECT 70.160 -81.120 71.400 -80.950 ;
        RECT 70.160 -81.350 70.330 -81.120 ;
        RECT 71.570 -81.290 71.740 -72.710 ;
        RECT 72.090 -80.710 72.260 -72.710 ;
        RECT 72.530 -80.710 72.700 -72.710 ;
        RECT 73.890 -73.040 74.060 -72.730 ;
        RECT 73.540 -73.210 74.060 -73.040 ;
        RECT 73.540 -76.150 73.710 -73.210 ;
        RECT 80.020 -76.120 80.190 -75.790 ;
        RECT 73.100 -80.260 73.270 -76.270 ;
        RECT 73.890 -78.270 74.060 -76.270 ;
        RECT 79.630 -78.250 79.800 -76.250 ;
        RECT 73.540 -80.260 73.710 -79.710 ;
        RECT 79.980 -80.260 80.150 -79.710 ;
        RECT 80.420 -80.260 80.590 -73.710 ;
        RECT 73.490 -80.760 73.660 -80.430 ;
        RECT 80.030 -80.770 80.200 -80.440 ;
        RECT 81.020 -80.710 81.190 -72.710 ;
        RECT 81.460 -80.710 81.630 -72.710 ;
        RECT 72.320 -81.090 72.650 -80.920 ;
        RECT 81.070 -81.080 81.400 -80.910 ;
        RECT 81.980 -80.950 82.150 -72.710 ;
        RECT 82.420 -80.710 82.590 -72.710 ;
        RECT 82.950 -80.710 83.120 -72.710 ;
        RECT 58.690 -81.460 61.450 -81.350 ;
        RECT 50.060 -83.880 50.230 -83.470 ;
        RECT 56.780 -85.700 56.950 -81.520 ;
        RECT 57.220 -81.960 57.390 -81.700 ;
        RECT 57.220 -82.130 57.430 -81.960 ;
        RECT 57.220 -83.580 57.390 -82.130 ;
        RECT 57.220 -83.750 57.430 -83.580 ;
        RECT 57.220 -85.700 57.390 -83.750 ;
        RECT 58.340 -85.700 58.510 -81.520 ;
        RECT 59.750 -81.520 61.450 -81.460 ;
        RECT 58.780 -81.970 58.950 -81.700 ;
        RECT 59.310 -81.970 59.480 -81.700 ;
        RECT 58.780 -82.140 58.970 -81.970 ;
        RECT 59.290 -82.140 59.480 -81.970 ;
        RECT 58.780 -83.590 58.950 -82.140 ;
        RECT 59.310 -83.590 59.480 -82.140 ;
        RECT 58.780 -83.760 59.480 -83.590 ;
        RECT 58.780 -85.700 58.950 -83.760 ;
        RECT 59.310 -85.700 59.480 -83.760 ;
        RECT 59.750 -85.700 59.920 -81.520 ;
        RECT 60.840 -81.960 61.010 -81.700 ;
        RECT 60.800 -82.130 61.010 -81.960 ;
        RECT 60.840 -83.610 61.010 -82.130 ;
        RECT 60.800 -83.780 61.010 -83.610 ;
        RECT 60.840 -85.700 61.010 -83.780 ;
        RECT 61.280 -85.700 61.450 -81.520 ;
        RECT 68.600 -81.520 70.330 -81.350 ;
        RECT 70.510 -81.350 71.740 -81.290 ;
        RECT 81.980 -81.120 83.220 -80.950 ;
        RECT 81.980 -81.350 82.150 -81.120 ;
        RECT 83.390 -81.290 83.560 -72.710 ;
        RECT 83.910 -80.710 84.080 -72.710 ;
        RECT 84.350 -80.710 84.520 -72.710 ;
        RECT 85.710 -73.040 85.880 -72.730 ;
        RECT 85.360 -73.210 85.880 -73.040 ;
        RECT 85.360 -76.150 85.530 -73.210 ;
        RECT 91.860 -76.120 92.030 -75.790 ;
        RECT 84.920 -80.260 85.090 -76.270 ;
        RECT 85.710 -78.270 85.880 -76.270 ;
        RECT 91.470 -78.250 91.640 -76.250 ;
        RECT 85.360 -80.260 85.530 -79.710 ;
        RECT 91.820 -80.260 91.990 -79.710 ;
        RECT 92.260 -80.260 92.430 -73.710 ;
        RECT 85.310 -80.760 85.480 -80.430 ;
        RECT 91.870 -80.770 92.040 -80.440 ;
        RECT 92.860 -80.710 93.030 -72.710 ;
        RECT 93.300 -80.710 93.470 -72.710 ;
        RECT 84.140 -81.090 84.470 -80.920 ;
        RECT 92.910 -81.080 93.240 -80.910 ;
        RECT 93.820 -80.950 93.990 -72.710 ;
        RECT 94.260 -80.710 94.430 -72.710 ;
        RECT 94.790 -80.710 94.960 -72.710 ;
        RECT 70.510 -81.460 73.270 -81.350 ;
        RECT 61.880 -83.880 62.050 -83.470 ;
        RECT 68.600 -85.700 68.770 -81.520 ;
        RECT 69.040 -81.960 69.210 -81.700 ;
        RECT 69.040 -82.130 69.250 -81.960 ;
        RECT 69.040 -83.580 69.210 -82.130 ;
        RECT 69.040 -83.750 69.250 -83.580 ;
        RECT 69.040 -85.700 69.210 -83.750 ;
        RECT 70.160 -85.700 70.330 -81.520 ;
        RECT 71.570 -81.520 73.270 -81.460 ;
        RECT 70.600 -81.970 70.770 -81.700 ;
        RECT 71.130 -81.970 71.300 -81.700 ;
        RECT 70.600 -82.140 70.790 -81.970 ;
        RECT 71.110 -82.140 71.300 -81.970 ;
        RECT 70.600 -83.590 70.770 -82.140 ;
        RECT 71.130 -83.590 71.300 -82.140 ;
        RECT 70.600 -83.760 71.300 -83.590 ;
        RECT 70.600 -85.700 70.770 -83.760 ;
        RECT 71.130 -85.700 71.300 -83.760 ;
        RECT 71.570 -85.700 71.740 -81.520 ;
        RECT 72.660 -81.960 72.830 -81.700 ;
        RECT 72.620 -82.130 72.830 -81.960 ;
        RECT 72.660 -83.610 72.830 -82.130 ;
        RECT 72.620 -83.780 72.830 -83.610 ;
        RECT 72.660 -85.700 72.830 -83.780 ;
        RECT 73.100 -85.700 73.270 -81.520 ;
        RECT 80.420 -81.520 82.150 -81.350 ;
        RECT 82.330 -81.350 83.560 -81.290 ;
        RECT 93.820 -81.120 95.060 -80.950 ;
        RECT 93.820 -81.350 93.990 -81.120 ;
        RECT 95.230 -81.290 95.400 -72.710 ;
        RECT 95.750 -80.710 95.920 -72.710 ;
        RECT 96.190 -80.710 96.360 -72.710 ;
        RECT 97.550 -73.040 97.720 -72.730 ;
        RECT 97.200 -73.210 97.720 -73.040 ;
        RECT 97.200 -76.150 97.370 -73.210 ;
        RECT 103.700 -76.120 103.870 -75.790 ;
        RECT 96.760 -80.260 96.930 -76.270 ;
        RECT 97.550 -78.270 97.720 -76.270 ;
        RECT 103.310 -78.250 103.480 -76.250 ;
        RECT 97.200 -80.260 97.370 -79.710 ;
        RECT 103.660 -80.260 103.830 -79.710 ;
        RECT 104.100 -80.260 104.270 -73.710 ;
        RECT 97.150 -80.760 97.320 -80.430 ;
        RECT 103.710 -80.770 103.880 -80.440 ;
        RECT 104.700 -80.710 104.870 -72.710 ;
        RECT 105.140 -80.710 105.310 -72.710 ;
        RECT 95.980 -81.090 96.310 -80.920 ;
        RECT 104.750 -81.080 105.080 -80.910 ;
        RECT 105.660 -80.950 105.830 -72.710 ;
        RECT 106.100 -80.710 106.270 -72.710 ;
        RECT 106.630 -80.710 106.800 -72.710 ;
        RECT 82.330 -81.460 85.090 -81.350 ;
        RECT 73.700 -83.880 73.870 -83.470 ;
        RECT 80.420 -85.700 80.590 -81.520 ;
        RECT 80.860 -81.960 81.030 -81.700 ;
        RECT 80.860 -82.130 81.070 -81.960 ;
        RECT 80.860 -83.580 81.030 -82.130 ;
        RECT 80.860 -83.750 81.070 -83.580 ;
        RECT 80.860 -85.700 81.030 -83.750 ;
        RECT 81.980 -85.700 82.150 -81.520 ;
        RECT 83.390 -81.520 85.090 -81.460 ;
        RECT 82.420 -81.970 82.590 -81.700 ;
        RECT 82.950 -81.970 83.120 -81.700 ;
        RECT 82.420 -82.140 82.610 -81.970 ;
        RECT 82.930 -82.140 83.120 -81.970 ;
        RECT 82.420 -83.590 82.590 -82.140 ;
        RECT 82.950 -83.590 83.120 -82.140 ;
        RECT 82.420 -83.760 83.120 -83.590 ;
        RECT 82.420 -85.700 82.590 -83.760 ;
        RECT 82.950 -85.700 83.120 -83.760 ;
        RECT 83.390 -85.700 83.560 -81.520 ;
        RECT 84.480 -81.960 84.650 -81.700 ;
        RECT 84.440 -82.130 84.650 -81.960 ;
        RECT 84.480 -83.610 84.650 -82.130 ;
        RECT 84.440 -83.780 84.650 -83.610 ;
        RECT 84.480 -85.700 84.650 -83.780 ;
        RECT 84.920 -85.700 85.090 -81.520 ;
        RECT 92.260 -81.520 93.990 -81.350 ;
        RECT 94.170 -81.350 95.400 -81.290 ;
        RECT 105.660 -81.120 106.900 -80.950 ;
        RECT 105.660 -81.350 105.830 -81.120 ;
        RECT 107.070 -81.290 107.240 -72.710 ;
        RECT 107.590 -80.710 107.760 -72.710 ;
        RECT 108.030 -80.710 108.200 -72.710 ;
        RECT 109.390 -73.040 109.560 -72.730 ;
        RECT 109.040 -73.210 109.560 -73.040 ;
        RECT 109.040 -76.150 109.210 -73.210 ;
        RECT 115.570 -76.120 115.740 -75.790 ;
        RECT 108.600 -80.260 108.770 -76.270 ;
        RECT 109.390 -78.270 109.560 -76.270 ;
        RECT 115.180 -78.250 115.350 -76.250 ;
        RECT 109.040 -80.260 109.210 -79.710 ;
        RECT 115.530 -80.260 115.700 -79.710 ;
        RECT 115.970 -80.260 116.140 -73.710 ;
        RECT 108.990 -80.760 109.160 -80.430 ;
        RECT 115.580 -80.770 115.750 -80.440 ;
        RECT 116.570 -80.710 116.740 -72.710 ;
        RECT 117.010 -80.710 117.180 -72.710 ;
        RECT 107.820 -81.090 108.150 -80.920 ;
        RECT 116.620 -81.080 116.950 -80.910 ;
        RECT 117.530 -80.950 117.700 -72.710 ;
        RECT 117.970 -80.710 118.140 -72.710 ;
        RECT 118.500 -80.710 118.670 -72.710 ;
        RECT 94.170 -81.460 96.930 -81.350 ;
        RECT 85.520 -83.880 85.690 -83.470 ;
        RECT 92.260 -85.700 92.430 -81.520 ;
        RECT 92.700 -81.960 92.870 -81.700 ;
        RECT 92.700 -82.130 92.910 -81.960 ;
        RECT 92.700 -83.580 92.870 -82.130 ;
        RECT 92.700 -83.750 92.910 -83.580 ;
        RECT 92.700 -85.700 92.870 -83.750 ;
        RECT 93.820 -85.700 93.990 -81.520 ;
        RECT 95.230 -81.520 96.930 -81.460 ;
        RECT 94.260 -81.970 94.430 -81.700 ;
        RECT 94.790 -81.970 94.960 -81.700 ;
        RECT 94.260 -82.140 94.450 -81.970 ;
        RECT 94.770 -82.140 94.960 -81.970 ;
        RECT 94.260 -83.590 94.430 -82.140 ;
        RECT 94.790 -83.590 94.960 -82.140 ;
        RECT 94.260 -83.760 94.960 -83.590 ;
        RECT 94.260 -85.700 94.430 -83.760 ;
        RECT 94.790 -85.700 94.960 -83.760 ;
        RECT 95.230 -85.700 95.400 -81.520 ;
        RECT 96.320 -81.960 96.490 -81.700 ;
        RECT 96.280 -82.130 96.490 -81.960 ;
        RECT 96.320 -83.610 96.490 -82.130 ;
        RECT 96.280 -83.780 96.490 -83.610 ;
        RECT 96.320 -85.700 96.490 -83.780 ;
        RECT 96.760 -85.700 96.930 -81.520 ;
        RECT 104.100 -81.520 105.830 -81.350 ;
        RECT 106.010 -81.350 107.240 -81.290 ;
        RECT 117.530 -81.120 118.770 -80.950 ;
        RECT 117.530 -81.350 117.700 -81.120 ;
        RECT 118.940 -81.290 119.110 -72.710 ;
        RECT 119.460 -80.710 119.630 -72.710 ;
        RECT 119.900 -80.710 120.070 -72.710 ;
        RECT 121.260 -73.040 121.430 -72.730 ;
        RECT 120.910 -73.210 121.430 -73.040 ;
        RECT 120.910 -76.150 121.080 -73.210 ;
        RECT 127.440 -76.120 127.610 -75.790 ;
        RECT 120.470 -80.260 120.640 -76.270 ;
        RECT 121.260 -78.270 121.430 -76.270 ;
        RECT 127.050 -78.250 127.220 -76.250 ;
        RECT 120.910 -80.260 121.080 -79.710 ;
        RECT 127.400 -80.260 127.570 -79.710 ;
        RECT 127.840 -80.260 128.010 -73.710 ;
        RECT 120.860 -80.760 121.030 -80.430 ;
        RECT 127.450 -80.770 127.620 -80.440 ;
        RECT 128.440 -80.710 128.610 -72.710 ;
        RECT 128.880 -80.710 129.050 -72.710 ;
        RECT 119.690 -81.090 120.020 -80.920 ;
        RECT 128.490 -81.080 128.820 -80.910 ;
        RECT 129.400 -80.950 129.570 -72.710 ;
        RECT 129.840 -80.710 130.010 -72.710 ;
        RECT 130.370 -80.710 130.540 -72.710 ;
        RECT 106.010 -81.460 108.770 -81.350 ;
        RECT 97.360 -83.880 97.530 -83.470 ;
        RECT 104.100 -85.700 104.270 -81.520 ;
        RECT 104.540 -81.960 104.710 -81.700 ;
        RECT 104.540 -82.130 104.750 -81.960 ;
        RECT 104.540 -83.580 104.710 -82.130 ;
        RECT 104.540 -83.750 104.750 -83.580 ;
        RECT 104.540 -85.700 104.710 -83.750 ;
        RECT 105.660 -85.700 105.830 -81.520 ;
        RECT 107.070 -81.520 108.770 -81.460 ;
        RECT 106.100 -81.970 106.270 -81.700 ;
        RECT 106.630 -81.970 106.800 -81.700 ;
        RECT 106.100 -82.140 106.290 -81.970 ;
        RECT 106.610 -82.140 106.800 -81.970 ;
        RECT 106.100 -83.590 106.270 -82.140 ;
        RECT 106.630 -83.590 106.800 -82.140 ;
        RECT 106.100 -83.760 106.800 -83.590 ;
        RECT 106.100 -85.700 106.270 -83.760 ;
        RECT 106.630 -85.700 106.800 -83.760 ;
        RECT 107.070 -85.700 107.240 -81.520 ;
        RECT 108.160 -81.960 108.330 -81.700 ;
        RECT 108.120 -82.130 108.330 -81.960 ;
        RECT 108.160 -83.610 108.330 -82.130 ;
        RECT 108.120 -83.780 108.330 -83.610 ;
        RECT 108.160 -85.700 108.330 -83.780 ;
        RECT 108.600 -85.700 108.770 -81.520 ;
        RECT 115.970 -81.520 117.700 -81.350 ;
        RECT 117.880 -81.350 119.110 -81.290 ;
        RECT 129.400 -81.120 130.640 -80.950 ;
        RECT 129.400 -81.350 129.570 -81.120 ;
        RECT 130.810 -81.290 130.980 -72.710 ;
        RECT 131.330 -80.710 131.500 -72.710 ;
        RECT 131.770 -80.710 131.940 -72.710 ;
        RECT 133.130 -73.040 133.300 -72.730 ;
        RECT 132.780 -73.210 133.300 -73.040 ;
        RECT 132.780 -76.150 132.950 -73.210 ;
        RECT 136.450 -76.120 136.620 -75.790 ;
        RECT 132.340 -80.260 132.510 -76.270 ;
        RECT 133.130 -78.270 133.300 -76.270 ;
        RECT 136.060 -78.250 136.230 -76.250 ;
        RECT 132.780 -80.260 132.950 -79.710 ;
        RECT 136.410 -80.260 136.580 -79.710 ;
        RECT 136.850 -80.260 137.020 -73.710 ;
        RECT 132.730 -80.760 132.900 -80.430 ;
        RECT 136.460 -80.770 136.630 -80.440 ;
        RECT 137.450 -80.710 137.620 -72.710 ;
        RECT 137.890 -80.710 138.060 -72.710 ;
        RECT 131.560 -81.090 131.890 -80.920 ;
        RECT 137.500 -81.080 137.830 -80.910 ;
        RECT 138.410 -80.950 138.580 -72.710 ;
        RECT 138.850 -80.710 139.020 -72.710 ;
        RECT 139.380 -80.710 139.550 -72.710 ;
        RECT 117.880 -81.460 120.640 -81.350 ;
        RECT 109.200 -83.880 109.370 -83.470 ;
        RECT 115.970 -85.700 116.140 -81.520 ;
        RECT 116.410 -81.960 116.580 -81.700 ;
        RECT 116.410 -82.130 116.620 -81.960 ;
        RECT 116.410 -83.580 116.580 -82.130 ;
        RECT 116.410 -83.750 116.620 -83.580 ;
        RECT 116.410 -85.700 116.580 -83.750 ;
        RECT 117.530 -85.700 117.700 -81.520 ;
        RECT 118.940 -81.520 120.640 -81.460 ;
        RECT 117.970 -81.970 118.140 -81.700 ;
        RECT 118.500 -81.970 118.670 -81.700 ;
        RECT 117.970 -82.140 118.160 -81.970 ;
        RECT 118.480 -82.140 118.670 -81.970 ;
        RECT 117.970 -83.590 118.140 -82.140 ;
        RECT 118.500 -83.590 118.670 -82.140 ;
        RECT 117.970 -83.760 118.670 -83.590 ;
        RECT 117.970 -85.700 118.140 -83.760 ;
        RECT 118.500 -85.700 118.670 -83.760 ;
        RECT 118.940 -85.700 119.110 -81.520 ;
        RECT 120.030 -81.960 120.200 -81.700 ;
        RECT 119.990 -82.130 120.200 -81.960 ;
        RECT 120.030 -83.610 120.200 -82.130 ;
        RECT 119.990 -83.780 120.200 -83.610 ;
        RECT 120.030 -85.700 120.200 -83.780 ;
        RECT 120.470 -85.700 120.640 -81.520 ;
        RECT 127.840 -81.520 129.570 -81.350 ;
        RECT 129.750 -81.350 130.980 -81.290 ;
        RECT 138.410 -81.120 139.650 -80.950 ;
        RECT 138.410 -81.350 138.580 -81.120 ;
        RECT 139.820 -81.290 139.990 -72.710 ;
        RECT 140.340 -80.710 140.510 -72.710 ;
        RECT 140.780 -80.710 140.950 -72.710 ;
        RECT 142.140 -73.040 142.310 -72.730 ;
        RECT 141.790 -73.210 142.310 -73.040 ;
        RECT 141.790 -76.150 141.960 -73.210 ;
        RECT 141.350 -80.260 141.520 -76.270 ;
        RECT 142.140 -78.270 142.310 -76.270 ;
        RECT 141.790 -80.260 141.960 -79.710 ;
        RECT 141.740 -80.760 141.910 -80.430 ;
        RECT 140.570 -81.090 140.900 -80.920 ;
        RECT 129.750 -81.460 132.510 -81.350 ;
        RECT 121.070 -83.880 121.240 -83.470 ;
        RECT 127.840 -85.700 128.010 -81.520 ;
        RECT 128.280 -81.960 128.450 -81.700 ;
        RECT 128.280 -82.130 128.490 -81.960 ;
        RECT 128.280 -83.580 128.450 -82.130 ;
        RECT 128.280 -83.750 128.490 -83.580 ;
        RECT 128.280 -85.700 128.450 -83.750 ;
        RECT 129.400 -85.700 129.570 -81.520 ;
        RECT 130.810 -81.520 132.510 -81.460 ;
        RECT 129.840 -81.970 130.010 -81.700 ;
        RECT 130.370 -81.970 130.540 -81.700 ;
        RECT 129.840 -82.140 130.030 -81.970 ;
        RECT 130.350 -82.140 130.540 -81.970 ;
        RECT 129.840 -83.590 130.010 -82.140 ;
        RECT 130.370 -83.590 130.540 -82.140 ;
        RECT 129.840 -83.760 130.540 -83.590 ;
        RECT 129.840 -85.700 130.010 -83.760 ;
        RECT 130.370 -85.700 130.540 -83.760 ;
        RECT 130.810 -85.700 130.980 -81.520 ;
        RECT 131.900 -81.960 132.070 -81.700 ;
        RECT 131.860 -82.130 132.070 -81.960 ;
        RECT 131.900 -83.610 132.070 -82.130 ;
        RECT 131.860 -83.780 132.070 -83.610 ;
        RECT 131.900 -85.700 132.070 -83.780 ;
        RECT 132.340 -85.700 132.510 -81.520 ;
        RECT 136.850 -81.520 138.580 -81.350 ;
        RECT 138.760 -81.350 139.990 -81.290 ;
        RECT 138.760 -81.460 141.520 -81.350 ;
        RECT 132.940 -83.880 133.110 -83.470 ;
        RECT 136.850 -85.700 137.020 -81.520 ;
        RECT 137.290 -81.960 137.460 -81.700 ;
        RECT 137.290 -82.130 137.500 -81.960 ;
        RECT 137.290 -83.580 137.460 -82.130 ;
        RECT 137.290 -83.750 137.500 -83.580 ;
        RECT 137.290 -85.700 137.460 -83.750 ;
        RECT 138.410 -85.700 138.580 -81.520 ;
        RECT 139.820 -81.520 141.520 -81.460 ;
        RECT 138.850 -81.970 139.020 -81.700 ;
        RECT 139.380 -81.970 139.550 -81.700 ;
        RECT 138.850 -82.140 139.040 -81.970 ;
        RECT 139.360 -82.140 139.550 -81.970 ;
        RECT 138.850 -83.590 139.020 -82.140 ;
        RECT 139.380 -83.590 139.550 -82.140 ;
        RECT 138.850 -83.760 139.550 -83.590 ;
        RECT 138.850 -85.700 139.020 -83.760 ;
        RECT 139.380 -85.700 139.550 -83.760 ;
        RECT 139.820 -85.700 139.990 -81.520 ;
        RECT 140.910 -81.960 141.080 -81.700 ;
        RECT 140.870 -82.130 141.080 -81.960 ;
        RECT 140.910 -83.610 141.080 -82.130 ;
        RECT 140.870 -83.780 141.080 -83.610 ;
        RECT 140.910 -85.700 141.080 -83.780 ;
        RECT 141.350 -85.700 141.520 -81.520 ;
        RECT 141.950 -83.880 142.120 -83.470 ;
        RECT -37.290 -86.120 -36.960 -85.950 ;
        RECT -33.240 -86.120 -32.910 -85.950 ;
        RECT -25.790 -86.120 -25.460 -85.950 ;
        RECT -21.740 -86.120 -21.410 -85.950 ;
        RECT -13.970 -86.120 -13.640 -85.950 ;
        RECT -9.920 -86.120 -9.590 -85.950 ;
        RECT -2.160 -86.120 -1.830 -85.950 ;
        RECT 1.890 -86.120 2.220 -85.950 ;
        RECT 9.650 -86.120 9.980 -85.950 ;
        RECT 13.700 -86.120 14.030 -85.950 ;
        RECT 21.470 -86.120 21.800 -85.950 ;
        RECT 25.520 -86.120 25.850 -85.950 ;
        RECT 33.290 -86.120 33.620 -85.950 ;
        RECT 37.340 -86.120 37.670 -85.950 ;
        RECT 45.110 -86.120 45.440 -85.950 ;
        RECT 49.160 -86.120 49.490 -85.950 ;
        RECT 56.930 -86.120 57.260 -85.950 ;
        RECT 60.980 -86.120 61.310 -85.950 ;
        RECT 68.750 -86.120 69.080 -85.950 ;
        RECT 72.800 -86.120 73.130 -85.950 ;
        RECT 80.570 -86.120 80.900 -85.950 ;
        RECT 84.620 -86.120 84.950 -85.950 ;
        RECT 92.410 -86.120 92.740 -85.950 ;
        RECT 96.460 -86.120 96.790 -85.950 ;
        RECT 104.250 -86.120 104.580 -85.950 ;
        RECT 108.300 -86.120 108.630 -85.950 ;
        RECT 116.120 -86.120 116.450 -85.950 ;
        RECT 120.170 -86.120 120.500 -85.950 ;
        RECT 127.990 -86.120 128.320 -85.950 ;
        RECT 132.040 -86.120 132.370 -85.950 ;
        RECT 137.000 -86.120 137.330 -85.950 ;
        RECT 141.050 -86.120 141.380 -85.950 ;
      LAYER mcon ;
        RECT 4.420 49.990 4.590 50.160 ;
        RECT 5.290 49.990 5.460 50.160 ;
        RECT 6.160 49.990 6.330 50.160 ;
        RECT 10.170 49.990 10.340 50.160 ;
        RECT 11.040 49.990 11.210 50.160 ;
        RECT 11.910 49.990 12.080 50.160 ;
        RECT 15.920 49.990 16.090 50.160 ;
        RECT 16.790 49.990 16.960 50.160 ;
        RECT 17.660 49.990 17.830 50.160 ;
        RECT 21.670 49.990 21.840 50.160 ;
        RECT 22.540 49.990 22.710 50.160 ;
        RECT 23.410 49.990 23.580 50.160 ;
        RECT 27.420 49.990 27.590 50.160 ;
        RECT 28.290 49.990 28.460 50.160 ;
        RECT 29.160 49.990 29.330 50.160 ;
        RECT 33.170 49.990 33.340 50.160 ;
        RECT 34.040 49.990 34.210 50.160 ;
        RECT 34.910 49.990 35.080 50.160 ;
        RECT 38.920 49.990 39.090 50.160 ;
        RECT 39.790 49.990 39.960 50.160 ;
        RECT 40.660 49.990 40.830 50.160 ;
        RECT 44.670 49.990 44.840 50.160 ;
        RECT 45.540 49.990 45.710 50.160 ;
        RECT 46.410 49.990 46.580 50.160 ;
        RECT 50.420 49.990 50.590 50.160 ;
        RECT 51.290 49.990 51.460 50.160 ;
        RECT 52.160 49.990 52.330 50.160 ;
        RECT 56.170 49.990 56.340 50.160 ;
        RECT 57.040 49.990 57.210 50.160 ;
        RECT 57.910 49.990 58.080 50.160 ;
        RECT 61.920 49.990 62.090 50.160 ;
        RECT 62.790 49.990 62.960 50.160 ;
        RECT 63.660 49.990 63.830 50.160 ;
        RECT 67.670 49.990 67.840 50.160 ;
        RECT 68.540 49.990 68.710 50.160 ;
        RECT 69.410 49.990 69.580 50.160 ;
        RECT 73.420 49.990 73.590 50.160 ;
        RECT 74.290 49.990 74.460 50.160 ;
        RECT 75.160 49.990 75.330 50.160 ;
        RECT 79.170 49.990 79.340 50.160 ;
        RECT 80.040 49.990 80.210 50.160 ;
        RECT 80.910 49.990 81.080 50.160 ;
        RECT 84.920 49.990 85.090 50.160 ;
        RECT 85.790 49.990 85.960 50.160 ;
        RECT 86.660 49.990 86.830 50.160 ;
        RECT 90.670 49.990 90.840 50.160 ;
        RECT 91.540 49.990 91.710 50.160 ;
        RECT 92.410 49.990 92.580 50.160 ;
        RECT 4.110 49.460 4.280 49.630 ;
        RECT 5.320 49.480 5.490 49.650 ;
        RECT 6.470 49.460 6.640 49.630 ;
        RECT 9.860 49.460 10.030 49.630 ;
        RECT 11.070 49.480 11.240 49.650 ;
        RECT 12.220 49.460 12.390 49.630 ;
        RECT 15.610 49.460 15.780 49.630 ;
        RECT 16.820 49.480 16.990 49.650 ;
        RECT 17.970 49.460 18.140 49.630 ;
        RECT 21.360 49.460 21.530 49.630 ;
        RECT 22.570 49.480 22.740 49.650 ;
        RECT 23.720 49.460 23.890 49.630 ;
        RECT 27.110 49.460 27.280 49.630 ;
        RECT 28.320 49.480 28.490 49.650 ;
        RECT 29.470 49.460 29.640 49.630 ;
        RECT 32.860 49.460 33.030 49.630 ;
        RECT 34.070 49.480 34.240 49.650 ;
        RECT 35.220 49.460 35.390 49.630 ;
        RECT 38.610 49.460 38.780 49.630 ;
        RECT 39.820 49.480 39.990 49.650 ;
        RECT 40.970 49.460 41.140 49.630 ;
        RECT 44.360 49.460 44.530 49.630 ;
        RECT 45.570 49.480 45.740 49.650 ;
        RECT 46.720 49.460 46.890 49.630 ;
        RECT 50.110 49.460 50.280 49.630 ;
        RECT 51.320 49.480 51.490 49.650 ;
        RECT 52.470 49.460 52.640 49.630 ;
        RECT 55.860 49.460 56.030 49.630 ;
        RECT 57.070 49.480 57.240 49.650 ;
        RECT 58.220 49.460 58.390 49.630 ;
        RECT 61.610 49.460 61.780 49.630 ;
        RECT 62.820 49.480 62.990 49.650 ;
        RECT 63.970 49.460 64.140 49.630 ;
        RECT 67.360 49.460 67.530 49.630 ;
        RECT 68.570 49.480 68.740 49.650 ;
        RECT 69.720 49.460 69.890 49.630 ;
        RECT 73.110 49.460 73.280 49.630 ;
        RECT 74.320 49.480 74.490 49.650 ;
        RECT 75.470 49.460 75.640 49.630 ;
        RECT 78.860 49.460 79.030 49.630 ;
        RECT 80.070 49.480 80.240 49.650 ;
        RECT 81.220 49.460 81.390 49.630 ;
        RECT 84.610 49.460 84.780 49.630 ;
        RECT 85.820 49.480 85.990 49.650 ;
        RECT 86.970 49.460 87.140 49.630 ;
        RECT 90.360 49.460 90.530 49.630 ;
        RECT 91.570 49.480 91.740 49.650 ;
        RECT 92.720 49.460 92.890 49.630 ;
        RECT 7.120 48.250 7.290 48.420 ;
        RECT 3.030 48.050 3.200 48.220 ;
        RECT 3.950 48.050 4.120 48.220 ;
        RECT 5.580 47.960 5.750 48.130 ;
        RECT 12.870 48.250 13.040 48.420 ;
        RECT 2.520 47.610 2.690 47.780 ;
        RECT 8.780 48.050 8.950 48.220 ;
        RECT 9.700 48.050 9.870 48.220 ;
        RECT 11.330 47.960 11.500 48.130 ;
        RECT 18.620 48.250 18.790 48.420 ;
        RECT 8.270 47.610 8.440 47.780 ;
        RECT 3.420 46.420 3.590 46.590 ;
        RECT 6.110 47.130 6.280 47.300 ;
        RECT 14.530 48.050 14.700 48.220 ;
        RECT 15.450 48.050 15.620 48.220 ;
        RECT 17.080 47.960 17.250 48.130 ;
        RECT 24.370 48.250 24.540 48.420 ;
        RECT 14.020 47.610 14.190 47.780 ;
        RECT 8.060 46.790 8.230 46.960 ;
        RECT 5.010 46.380 5.180 46.550 ;
        RECT 6.650 46.380 6.820 46.550 ;
        RECT 7.560 46.380 7.730 46.550 ;
        RECT 9.170 46.420 9.340 46.590 ;
        RECT 11.860 47.130 12.030 47.300 ;
        RECT 20.280 48.050 20.450 48.220 ;
        RECT 21.200 48.050 21.370 48.220 ;
        RECT 22.830 47.960 23.000 48.130 ;
        RECT 30.120 48.250 30.290 48.420 ;
        RECT 19.770 47.610 19.940 47.780 ;
        RECT 13.810 46.790 13.980 46.960 ;
        RECT 10.760 46.380 10.930 46.550 ;
        RECT 12.400 46.380 12.570 46.550 ;
        RECT 13.310 46.380 13.480 46.550 ;
        RECT 14.920 46.420 15.090 46.590 ;
        RECT 17.610 47.130 17.780 47.300 ;
        RECT 26.030 48.050 26.200 48.220 ;
        RECT 26.950 48.050 27.120 48.220 ;
        RECT 28.580 47.960 28.750 48.130 ;
        RECT 35.870 48.250 36.040 48.420 ;
        RECT 25.520 47.610 25.690 47.780 ;
        RECT 19.560 46.790 19.730 46.960 ;
        RECT 16.510 46.380 16.680 46.550 ;
        RECT 18.150 46.380 18.320 46.550 ;
        RECT 19.060 46.380 19.230 46.550 ;
        RECT 20.670 46.420 20.840 46.590 ;
        RECT 23.360 47.130 23.530 47.300 ;
        RECT 31.780 48.050 31.950 48.220 ;
        RECT 32.700 48.050 32.870 48.220 ;
        RECT 34.330 47.960 34.500 48.130 ;
        RECT 41.620 48.250 41.790 48.420 ;
        RECT 31.270 47.610 31.440 47.780 ;
        RECT 25.310 46.790 25.480 46.960 ;
        RECT 22.260 46.380 22.430 46.550 ;
        RECT 23.900 46.380 24.070 46.550 ;
        RECT 24.810 46.380 24.980 46.550 ;
        RECT 26.420 46.420 26.590 46.590 ;
        RECT 29.110 47.130 29.280 47.300 ;
        RECT 37.530 48.050 37.700 48.220 ;
        RECT 38.450 48.050 38.620 48.220 ;
        RECT 40.080 47.960 40.250 48.130 ;
        RECT 47.370 48.250 47.540 48.420 ;
        RECT 37.020 47.610 37.190 47.780 ;
        RECT 31.060 46.790 31.230 46.960 ;
        RECT 28.010 46.380 28.180 46.550 ;
        RECT 29.650 46.380 29.820 46.550 ;
        RECT 30.560 46.380 30.730 46.550 ;
        RECT 32.170 46.420 32.340 46.590 ;
        RECT 34.860 47.130 35.030 47.300 ;
        RECT 43.280 48.050 43.450 48.220 ;
        RECT 44.200 48.050 44.370 48.220 ;
        RECT 45.830 47.960 46.000 48.130 ;
        RECT 53.120 48.250 53.290 48.420 ;
        RECT 42.770 47.610 42.940 47.780 ;
        RECT 36.810 46.790 36.980 46.960 ;
        RECT 33.760 46.380 33.930 46.550 ;
        RECT 35.400 46.380 35.570 46.550 ;
        RECT 36.310 46.380 36.480 46.550 ;
        RECT 37.920 46.420 38.090 46.590 ;
        RECT 40.610 47.130 40.780 47.300 ;
        RECT 49.030 48.050 49.200 48.220 ;
        RECT 49.950 48.050 50.120 48.220 ;
        RECT 51.580 47.960 51.750 48.130 ;
        RECT 58.870 48.250 59.040 48.420 ;
        RECT 48.520 47.610 48.690 47.780 ;
        RECT 42.560 46.790 42.730 46.960 ;
        RECT 39.510 46.380 39.680 46.550 ;
        RECT 41.150 46.380 41.320 46.550 ;
        RECT 42.060 46.380 42.230 46.550 ;
        RECT 43.670 46.420 43.840 46.590 ;
        RECT 46.360 47.130 46.530 47.300 ;
        RECT 54.780 48.050 54.950 48.220 ;
        RECT 55.700 48.050 55.870 48.220 ;
        RECT 57.330 47.960 57.500 48.130 ;
        RECT 64.620 48.250 64.790 48.420 ;
        RECT 54.270 47.610 54.440 47.780 ;
        RECT 48.310 46.790 48.480 46.960 ;
        RECT 45.260 46.380 45.430 46.550 ;
        RECT 46.900 46.380 47.070 46.550 ;
        RECT 47.810 46.380 47.980 46.550 ;
        RECT 49.420 46.420 49.590 46.590 ;
        RECT 52.110 47.130 52.280 47.300 ;
        RECT 60.530 48.050 60.700 48.220 ;
        RECT 61.450 48.050 61.620 48.220 ;
        RECT 63.080 47.960 63.250 48.130 ;
        RECT 70.370 48.250 70.540 48.420 ;
        RECT 60.020 47.610 60.190 47.780 ;
        RECT 54.060 46.790 54.230 46.960 ;
        RECT 51.010 46.380 51.180 46.550 ;
        RECT 52.650 46.380 52.820 46.550 ;
        RECT 53.560 46.380 53.730 46.550 ;
        RECT 55.170 46.420 55.340 46.590 ;
        RECT 57.860 47.130 58.030 47.300 ;
        RECT 66.280 48.050 66.450 48.220 ;
        RECT 67.200 48.050 67.370 48.220 ;
        RECT 68.830 47.960 69.000 48.130 ;
        RECT 76.120 48.250 76.290 48.420 ;
        RECT 65.770 47.610 65.940 47.780 ;
        RECT 59.810 46.790 59.980 46.960 ;
        RECT 56.760 46.380 56.930 46.550 ;
        RECT 58.400 46.380 58.570 46.550 ;
        RECT 59.310 46.380 59.480 46.550 ;
        RECT 60.920 46.420 61.090 46.590 ;
        RECT 63.610 47.130 63.780 47.300 ;
        RECT 72.030 48.050 72.200 48.220 ;
        RECT 72.950 48.050 73.120 48.220 ;
        RECT 74.580 47.960 74.750 48.130 ;
        RECT 81.870 48.250 82.040 48.420 ;
        RECT 71.520 47.610 71.690 47.780 ;
        RECT 65.560 46.790 65.730 46.960 ;
        RECT 62.510 46.380 62.680 46.550 ;
        RECT 64.150 46.380 64.320 46.550 ;
        RECT 65.060 46.380 65.230 46.550 ;
        RECT 66.670 46.420 66.840 46.590 ;
        RECT 69.360 47.130 69.530 47.300 ;
        RECT 77.780 48.050 77.950 48.220 ;
        RECT 78.700 48.050 78.870 48.220 ;
        RECT 80.330 47.960 80.500 48.130 ;
        RECT 87.620 48.250 87.790 48.420 ;
        RECT 77.270 47.610 77.440 47.780 ;
        RECT 71.310 46.790 71.480 46.960 ;
        RECT 68.260 46.380 68.430 46.550 ;
        RECT 69.900 46.380 70.070 46.550 ;
        RECT 70.810 46.380 70.980 46.550 ;
        RECT 72.420 46.420 72.590 46.590 ;
        RECT 75.110 47.130 75.280 47.300 ;
        RECT 83.530 48.050 83.700 48.220 ;
        RECT 84.450 48.050 84.620 48.220 ;
        RECT 86.080 47.960 86.250 48.130 ;
        RECT 93.370 48.250 93.540 48.420 ;
        RECT 83.020 47.610 83.190 47.780 ;
        RECT 77.060 46.790 77.230 46.960 ;
        RECT 74.010 46.380 74.180 46.550 ;
        RECT 75.650 46.380 75.820 46.550 ;
        RECT 76.560 46.380 76.730 46.550 ;
        RECT 78.170 46.420 78.340 46.590 ;
        RECT 80.860 47.130 81.030 47.300 ;
        RECT 89.280 48.050 89.450 48.220 ;
        RECT 90.200 48.050 90.370 48.220 ;
        RECT 91.830 47.960 92.000 48.130 ;
        RECT 88.770 47.610 88.940 47.780 ;
        RECT 82.810 46.790 82.980 46.960 ;
        RECT 79.760 46.380 79.930 46.550 ;
        RECT 81.400 46.380 81.570 46.550 ;
        RECT 82.310 46.380 82.480 46.550 ;
        RECT 83.920 46.420 84.090 46.590 ;
        RECT 86.610 47.130 86.780 47.300 ;
        RECT 88.560 46.790 88.730 46.960 ;
        RECT 85.510 46.380 85.680 46.550 ;
        RECT 87.150 46.380 87.320 46.550 ;
        RECT 88.060 46.380 88.230 46.550 ;
        RECT 89.670 46.420 89.840 46.590 ;
        RECT 92.360 47.130 92.530 47.300 ;
        RECT 94.310 46.790 94.480 46.960 ;
        RECT 91.260 46.380 91.430 46.550 ;
        RECT 92.900 46.380 93.070 46.550 ;
        RECT 93.810 46.380 93.980 46.550 ;
        RECT 7.120 45.840 7.290 46.010 ;
        RECT 3.030 45.640 3.200 45.810 ;
        RECT 3.950 45.640 4.120 45.810 ;
        RECT 5.580 45.550 5.750 45.720 ;
        RECT 12.870 45.840 13.040 46.010 ;
        RECT 2.520 45.200 2.690 45.370 ;
        RECT 8.780 45.640 8.950 45.810 ;
        RECT 9.700 45.640 9.870 45.810 ;
        RECT 11.330 45.550 11.500 45.720 ;
        RECT 18.620 45.840 18.790 46.010 ;
        RECT 8.270 45.200 8.440 45.370 ;
        RECT 3.420 44.010 3.590 44.180 ;
        RECT 6.110 44.720 6.280 44.890 ;
        RECT 14.530 45.640 14.700 45.810 ;
        RECT 15.450 45.640 15.620 45.810 ;
        RECT 17.080 45.550 17.250 45.720 ;
        RECT 24.370 45.840 24.540 46.010 ;
        RECT 14.020 45.200 14.190 45.370 ;
        RECT 8.060 44.380 8.230 44.550 ;
        RECT 5.010 43.970 5.180 44.140 ;
        RECT 6.650 43.970 6.820 44.140 ;
        RECT 7.560 43.970 7.730 44.140 ;
        RECT 7.120 43.110 7.290 43.280 ;
        RECT 9.170 44.010 9.340 44.180 ;
        RECT 11.860 44.720 12.030 44.890 ;
        RECT 20.280 45.640 20.450 45.810 ;
        RECT 21.200 45.640 21.370 45.810 ;
        RECT 22.830 45.550 23.000 45.720 ;
        RECT 30.120 45.840 30.290 46.010 ;
        RECT 19.770 45.200 19.940 45.370 ;
        RECT 13.810 44.380 13.980 44.550 ;
        RECT 10.760 43.970 10.930 44.140 ;
        RECT 12.400 43.970 12.570 44.140 ;
        RECT 13.310 43.970 13.480 44.140 ;
        RECT 3.030 42.670 3.200 42.840 ;
        RECT 3.950 42.670 4.120 42.840 ;
        RECT 5.580 42.580 5.750 42.750 ;
        RECT 12.870 43.110 13.040 43.280 ;
        RECT 14.920 44.010 15.090 44.180 ;
        RECT 17.610 44.720 17.780 44.890 ;
        RECT 26.030 45.640 26.200 45.810 ;
        RECT 26.950 45.640 27.120 45.810 ;
        RECT 28.580 45.550 28.750 45.720 ;
        RECT 35.870 45.840 36.040 46.010 ;
        RECT 25.520 45.200 25.690 45.370 ;
        RECT 19.560 44.380 19.730 44.550 ;
        RECT 16.510 43.970 16.680 44.140 ;
        RECT 18.150 43.970 18.320 44.140 ;
        RECT 19.060 43.970 19.230 44.140 ;
        RECT 2.520 42.230 2.690 42.400 ;
        RECT 8.780 42.670 8.950 42.840 ;
        RECT 9.700 42.670 9.870 42.840 ;
        RECT 11.330 42.580 11.500 42.750 ;
        RECT 18.620 43.110 18.790 43.280 ;
        RECT 20.670 44.010 20.840 44.180 ;
        RECT 23.360 44.720 23.530 44.890 ;
        RECT 31.780 45.640 31.950 45.810 ;
        RECT 32.700 45.640 32.870 45.810 ;
        RECT 34.330 45.550 34.500 45.720 ;
        RECT 41.620 45.840 41.790 46.010 ;
        RECT 31.270 45.200 31.440 45.370 ;
        RECT 25.310 44.380 25.480 44.550 ;
        RECT 22.260 43.970 22.430 44.140 ;
        RECT 23.900 43.970 24.070 44.140 ;
        RECT 24.810 43.970 24.980 44.140 ;
        RECT 8.270 42.230 8.440 42.400 ;
        RECT 3.420 41.040 3.590 41.210 ;
        RECT 6.110 41.750 6.280 41.920 ;
        RECT 14.530 42.670 14.700 42.840 ;
        RECT 15.450 42.670 15.620 42.840 ;
        RECT 17.080 42.580 17.250 42.750 ;
        RECT 24.370 43.110 24.540 43.280 ;
        RECT 26.420 44.010 26.590 44.180 ;
        RECT 29.110 44.720 29.280 44.890 ;
        RECT 37.530 45.640 37.700 45.810 ;
        RECT 38.450 45.640 38.620 45.810 ;
        RECT 40.080 45.550 40.250 45.720 ;
        RECT 47.370 45.840 47.540 46.010 ;
        RECT 37.020 45.200 37.190 45.370 ;
        RECT 31.060 44.380 31.230 44.550 ;
        RECT 28.010 43.970 28.180 44.140 ;
        RECT 29.650 43.970 29.820 44.140 ;
        RECT 30.560 43.970 30.730 44.140 ;
        RECT 14.020 42.230 14.190 42.400 ;
        RECT 8.060 41.410 8.230 41.580 ;
        RECT 5.010 41.000 5.180 41.170 ;
        RECT 6.650 41.000 6.820 41.170 ;
        RECT 7.560 41.000 7.730 41.170 ;
        RECT 9.170 41.040 9.340 41.210 ;
        RECT 11.860 41.750 12.030 41.920 ;
        RECT 20.280 42.670 20.450 42.840 ;
        RECT 21.200 42.670 21.370 42.840 ;
        RECT 22.830 42.580 23.000 42.750 ;
        RECT 30.120 43.110 30.290 43.280 ;
        RECT 32.170 44.010 32.340 44.180 ;
        RECT 34.860 44.720 35.030 44.890 ;
        RECT 43.280 45.640 43.450 45.810 ;
        RECT 44.200 45.640 44.370 45.810 ;
        RECT 45.830 45.550 46.000 45.720 ;
        RECT 53.120 45.840 53.290 46.010 ;
        RECT 42.770 45.200 42.940 45.370 ;
        RECT 36.810 44.380 36.980 44.550 ;
        RECT 33.760 43.970 33.930 44.140 ;
        RECT 35.400 43.970 35.570 44.140 ;
        RECT 36.310 43.970 36.480 44.140 ;
        RECT 19.770 42.230 19.940 42.400 ;
        RECT 13.810 41.410 13.980 41.580 ;
        RECT 10.760 41.000 10.930 41.170 ;
        RECT 12.400 41.000 12.570 41.170 ;
        RECT 13.310 41.000 13.480 41.170 ;
        RECT 14.920 41.040 15.090 41.210 ;
        RECT 17.610 41.750 17.780 41.920 ;
        RECT 26.030 42.670 26.200 42.840 ;
        RECT 26.950 42.670 27.120 42.840 ;
        RECT 28.580 42.580 28.750 42.750 ;
        RECT 35.870 43.110 36.040 43.280 ;
        RECT 37.920 44.010 38.090 44.180 ;
        RECT 40.610 44.720 40.780 44.890 ;
        RECT 49.030 45.640 49.200 45.810 ;
        RECT 49.950 45.640 50.120 45.810 ;
        RECT 51.580 45.550 51.750 45.720 ;
        RECT 58.870 45.840 59.040 46.010 ;
        RECT 48.520 45.200 48.690 45.370 ;
        RECT 42.560 44.380 42.730 44.550 ;
        RECT 39.510 43.970 39.680 44.140 ;
        RECT 41.150 43.970 41.320 44.140 ;
        RECT 42.060 43.970 42.230 44.140 ;
        RECT 25.520 42.230 25.690 42.400 ;
        RECT 19.560 41.410 19.730 41.580 ;
        RECT 16.510 41.000 16.680 41.170 ;
        RECT 18.150 41.000 18.320 41.170 ;
        RECT 19.060 41.000 19.230 41.170 ;
        RECT 20.670 41.040 20.840 41.210 ;
        RECT 23.360 41.750 23.530 41.920 ;
        RECT 31.780 42.670 31.950 42.840 ;
        RECT 32.700 42.670 32.870 42.840 ;
        RECT 34.330 42.580 34.500 42.750 ;
        RECT 41.620 43.110 41.790 43.280 ;
        RECT 43.670 44.010 43.840 44.180 ;
        RECT 46.360 44.720 46.530 44.890 ;
        RECT 54.780 45.640 54.950 45.810 ;
        RECT 55.700 45.640 55.870 45.810 ;
        RECT 57.330 45.550 57.500 45.720 ;
        RECT 64.620 45.840 64.790 46.010 ;
        RECT 54.270 45.200 54.440 45.370 ;
        RECT 48.310 44.380 48.480 44.550 ;
        RECT 45.260 43.970 45.430 44.140 ;
        RECT 46.900 43.970 47.070 44.140 ;
        RECT 47.810 43.970 47.980 44.140 ;
        RECT 31.270 42.230 31.440 42.400 ;
        RECT 25.310 41.410 25.480 41.580 ;
        RECT 22.260 41.000 22.430 41.170 ;
        RECT 23.900 41.000 24.070 41.170 ;
        RECT 24.810 41.000 24.980 41.170 ;
        RECT 26.420 41.040 26.590 41.210 ;
        RECT 29.110 41.750 29.280 41.920 ;
        RECT 37.530 42.670 37.700 42.840 ;
        RECT 38.450 42.670 38.620 42.840 ;
        RECT 40.080 42.580 40.250 42.750 ;
        RECT 47.370 43.110 47.540 43.280 ;
        RECT 49.420 44.010 49.590 44.180 ;
        RECT 52.110 44.720 52.280 44.890 ;
        RECT 60.530 45.640 60.700 45.810 ;
        RECT 61.450 45.640 61.620 45.810 ;
        RECT 63.080 45.550 63.250 45.720 ;
        RECT 70.370 45.840 70.540 46.010 ;
        RECT 60.020 45.200 60.190 45.370 ;
        RECT 54.060 44.380 54.230 44.550 ;
        RECT 51.010 43.970 51.180 44.140 ;
        RECT 52.650 43.970 52.820 44.140 ;
        RECT 53.560 43.970 53.730 44.140 ;
        RECT 37.020 42.230 37.190 42.400 ;
        RECT 31.060 41.410 31.230 41.580 ;
        RECT 28.010 41.000 28.180 41.170 ;
        RECT 29.650 41.000 29.820 41.170 ;
        RECT 30.560 41.000 30.730 41.170 ;
        RECT 32.170 41.040 32.340 41.210 ;
        RECT 34.860 41.750 35.030 41.920 ;
        RECT 43.280 42.670 43.450 42.840 ;
        RECT 44.200 42.670 44.370 42.840 ;
        RECT 45.830 42.580 46.000 42.750 ;
        RECT 53.120 43.110 53.290 43.280 ;
        RECT 55.170 44.010 55.340 44.180 ;
        RECT 57.860 44.720 58.030 44.890 ;
        RECT 66.280 45.640 66.450 45.810 ;
        RECT 67.200 45.640 67.370 45.810 ;
        RECT 68.830 45.550 69.000 45.720 ;
        RECT 76.120 45.840 76.290 46.010 ;
        RECT 65.770 45.200 65.940 45.370 ;
        RECT 59.810 44.380 59.980 44.550 ;
        RECT 56.760 43.970 56.930 44.140 ;
        RECT 58.400 43.970 58.570 44.140 ;
        RECT 59.310 43.970 59.480 44.140 ;
        RECT 42.770 42.230 42.940 42.400 ;
        RECT 36.810 41.410 36.980 41.580 ;
        RECT 33.760 41.000 33.930 41.170 ;
        RECT 35.400 41.000 35.570 41.170 ;
        RECT 36.310 41.000 36.480 41.170 ;
        RECT 37.920 41.040 38.090 41.210 ;
        RECT 40.610 41.750 40.780 41.920 ;
        RECT 49.030 42.670 49.200 42.840 ;
        RECT 49.950 42.670 50.120 42.840 ;
        RECT 51.580 42.580 51.750 42.750 ;
        RECT 58.870 43.110 59.040 43.280 ;
        RECT 60.920 44.010 61.090 44.180 ;
        RECT 63.610 44.720 63.780 44.890 ;
        RECT 72.030 45.640 72.200 45.810 ;
        RECT 72.950 45.640 73.120 45.810 ;
        RECT 74.580 45.550 74.750 45.720 ;
        RECT 81.870 45.840 82.040 46.010 ;
        RECT 71.520 45.200 71.690 45.370 ;
        RECT 65.560 44.380 65.730 44.550 ;
        RECT 62.510 43.970 62.680 44.140 ;
        RECT 64.150 43.970 64.320 44.140 ;
        RECT 65.060 43.970 65.230 44.140 ;
        RECT 48.520 42.230 48.690 42.400 ;
        RECT 42.560 41.410 42.730 41.580 ;
        RECT 39.510 41.000 39.680 41.170 ;
        RECT 41.150 41.000 41.320 41.170 ;
        RECT 42.060 41.000 42.230 41.170 ;
        RECT 43.670 41.040 43.840 41.210 ;
        RECT 46.360 41.750 46.530 41.920 ;
        RECT 54.780 42.670 54.950 42.840 ;
        RECT 55.700 42.670 55.870 42.840 ;
        RECT 57.330 42.580 57.500 42.750 ;
        RECT 64.620 43.110 64.790 43.280 ;
        RECT 66.670 44.010 66.840 44.180 ;
        RECT 69.360 44.720 69.530 44.890 ;
        RECT 77.780 45.640 77.950 45.810 ;
        RECT 78.700 45.640 78.870 45.810 ;
        RECT 80.330 45.550 80.500 45.720 ;
        RECT 87.620 45.840 87.790 46.010 ;
        RECT 77.270 45.200 77.440 45.370 ;
        RECT 71.310 44.380 71.480 44.550 ;
        RECT 68.260 43.970 68.430 44.140 ;
        RECT 69.900 43.970 70.070 44.140 ;
        RECT 70.810 43.970 70.980 44.140 ;
        RECT 54.270 42.230 54.440 42.400 ;
        RECT 48.310 41.410 48.480 41.580 ;
        RECT 45.260 41.000 45.430 41.170 ;
        RECT 46.900 41.000 47.070 41.170 ;
        RECT 47.810 41.000 47.980 41.170 ;
        RECT 49.420 41.040 49.590 41.210 ;
        RECT 52.110 41.750 52.280 41.920 ;
        RECT 60.530 42.670 60.700 42.840 ;
        RECT 61.450 42.670 61.620 42.840 ;
        RECT 63.080 42.580 63.250 42.750 ;
        RECT 70.370 43.110 70.540 43.280 ;
        RECT 72.420 44.010 72.590 44.180 ;
        RECT 75.110 44.720 75.280 44.890 ;
        RECT 83.530 45.640 83.700 45.810 ;
        RECT 84.450 45.640 84.620 45.810 ;
        RECT 86.080 45.550 86.250 45.720 ;
        RECT 93.370 45.840 93.540 46.010 ;
        RECT 83.020 45.200 83.190 45.370 ;
        RECT 77.060 44.380 77.230 44.550 ;
        RECT 74.010 43.970 74.180 44.140 ;
        RECT 75.650 43.970 75.820 44.140 ;
        RECT 76.560 43.970 76.730 44.140 ;
        RECT 60.020 42.230 60.190 42.400 ;
        RECT 54.060 41.410 54.230 41.580 ;
        RECT 51.010 41.000 51.180 41.170 ;
        RECT 52.650 41.000 52.820 41.170 ;
        RECT 53.560 41.000 53.730 41.170 ;
        RECT 55.170 41.040 55.340 41.210 ;
        RECT 57.860 41.750 58.030 41.920 ;
        RECT 66.280 42.670 66.450 42.840 ;
        RECT 67.200 42.670 67.370 42.840 ;
        RECT 68.830 42.580 69.000 42.750 ;
        RECT 76.120 43.110 76.290 43.280 ;
        RECT 78.170 44.010 78.340 44.180 ;
        RECT 80.860 44.720 81.030 44.890 ;
        RECT 89.280 45.640 89.450 45.810 ;
        RECT 90.200 45.640 90.370 45.810 ;
        RECT 91.830 45.550 92.000 45.720 ;
        RECT 88.770 45.200 88.940 45.370 ;
        RECT 82.810 44.380 82.980 44.550 ;
        RECT 79.760 43.970 79.930 44.140 ;
        RECT 81.400 43.970 81.570 44.140 ;
        RECT 82.310 43.970 82.480 44.140 ;
        RECT 65.770 42.230 65.940 42.400 ;
        RECT 59.810 41.410 59.980 41.580 ;
        RECT 56.760 41.000 56.930 41.170 ;
        RECT 58.400 41.000 58.570 41.170 ;
        RECT 59.310 41.000 59.480 41.170 ;
        RECT 60.920 41.040 61.090 41.210 ;
        RECT 63.610 41.750 63.780 41.920 ;
        RECT 72.030 42.670 72.200 42.840 ;
        RECT 72.950 42.670 73.120 42.840 ;
        RECT 74.580 42.580 74.750 42.750 ;
        RECT 81.870 43.110 82.040 43.280 ;
        RECT 83.920 44.010 84.090 44.180 ;
        RECT 86.610 44.720 86.780 44.890 ;
        RECT 88.560 44.380 88.730 44.550 ;
        RECT 85.510 43.970 85.680 44.140 ;
        RECT 87.150 43.970 87.320 44.140 ;
        RECT 88.060 43.970 88.230 44.140 ;
        RECT 71.520 42.230 71.690 42.400 ;
        RECT 65.560 41.410 65.730 41.580 ;
        RECT 62.510 41.000 62.680 41.170 ;
        RECT 64.150 41.000 64.320 41.170 ;
        RECT 65.060 41.000 65.230 41.170 ;
        RECT 66.670 41.040 66.840 41.210 ;
        RECT 69.360 41.750 69.530 41.920 ;
        RECT 77.780 42.670 77.950 42.840 ;
        RECT 78.700 42.670 78.870 42.840 ;
        RECT 80.330 42.580 80.500 42.750 ;
        RECT 87.620 43.110 87.790 43.280 ;
        RECT 89.670 44.010 89.840 44.180 ;
        RECT 92.360 44.720 92.530 44.890 ;
        RECT 94.310 44.380 94.480 44.550 ;
        RECT 91.260 43.970 91.430 44.140 ;
        RECT 92.900 43.970 93.070 44.140 ;
        RECT 93.810 43.970 93.980 44.140 ;
        RECT 77.270 42.230 77.440 42.400 ;
        RECT 71.310 41.410 71.480 41.580 ;
        RECT 68.260 41.000 68.430 41.170 ;
        RECT 69.900 41.000 70.070 41.170 ;
        RECT 70.810 41.000 70.980 41.170 ;
        RECT 72.420 41.040 72.590 41.210 ;
        RECT 75.110 41.750 75.280 41.920 ;
        RECT 83.530 42.670 83.700 42.840 ;
        RECT 84.450 42.670 84.620 42.840 ;
        RECT 86.080 42.580 86.250 42.750 ;
        RECT 83.020 42.230 83.190 42.400 ;
        RECT 77.060 41.410 77.230 41.580 ;
        RECT 74.010 41.000 74.180 41.170 ;
        RECT 75.650 41.000 75.820 41.170 ;
        RECT 76.560 41.000 76.730 41.170 ;
        RECT 78.170 41.040 78.340 41.210 ;
        RECT 80.860 41.750 81.030 41.920 ;
        RECT 89.280 42.670 89.450 42.840 ;
        RECT 90.200 42.670 90.370 42.840 ;
        RECT 91.830 42.580 92.000 42.750 ;
        RECT 88.770 42.230 88.940 42.400 ;
        RECT 82.810 41.410 82.980 41.580 ;
        RECT 79.760 41.000 79.930 41.170 ;
        RECT 81.400 41.000 81.570 41.170 ;
        RECT 82.310 41.000 82.480 41.170 ;
        RECT 83.920 41.040 84.090 41.210 ;
        RECT 86.610 41.750 86.780 41.920 ;
        RECT 88.560 41.410 88.730 41.580 ;
        RECT 85.510 41.000 85.680 41.170 ;
        RECT 87.150 41.000 87.320 41.170 ;
        RECT 88.060 41.000 88.230 41.170 ;
        RECT 89.670 41.040 89.840 41.210 ;
        RECT 92.360 41.750 92.530 41.920 ;
        RECT 94.310 41.410 94.480 41.580 ;
        RECT 91.260 41.000 91.430 41.170 ;
        RECT 92.900 41.000 93.070 41.170 ;
        RECT 93.810 41.000 93.980 41.170 ;
        RECT 7.120 40.460 7.290 40.630 ;
        RECT 3.030 40.260 3.200 40.430 ;
        RECT 3.950 40.260 4.120 40.430 ;
        RECT 5.580 40.170 5.750 40.340 ;
        RECT 12.870 40.460 13.040 40.630 ;
        RECT 2.520 39.820 2.690 39.990 ;
        RECT 8.780 40.260 8.950 40.430 ;
        RECT 9.700 40.260 9.870 40.430 ;
        RECT 11.330 40.170 11.500 40.340 ;
        RECT 18.620 40.460 18.790 40.630 ;
        RECT 8.270 39.820 8.440 39.990 ;
        RECT 3.420 38.630 3.590 38.800 ;
        RECT 6.110 39.340 6.280 39.510 ;
        RECT 14.530 40.260 14.700 40.430 ;
        RECT 15.450 40.260 15.620 40.430 ;
        RECT 17.080 40.170 17.250 40.340 ;
        RECT 24.370 40.460 24.540 40.630 ;
        RECT 14.020 39.820 14.190 39.990 ;
        RECT 8.060 39.000 8.230 39.170 ;
        RECT 5.010 38.590 5.180 38.760 ;
        RECT 6.650 38.590 6.820 38.760 ;
        RECT 7.560 38.590 7.730 38.760 ;
        RECT 9.170 38.630 9.340 38.800 ;
        RECT 11.860 39.340 12.030 39.510 ;
        RECT 20.280 40.260 20.450 40.430 ;
        RECT 21.200 40.260 21.370 40.430 ;
        RECT 22.830 40.170 23.000 40.340 ;
        RECT 30.120 40.460 30.290 40.630 ;
        RECT 19.770 39.820 19.940 39.990 ;
        RECT 13.810 39.000 13.980 39.170 ;
        RECT 10.760 38.590 10.930 38.760 ;
        RECT 12.400 38.590 12.570 38.760 ;
        RECT 13.310 38.590 13.480 38.760 ;
        RECT 14.920 38.630 15.090 38.800 ;
        RECT 17.610 39.340 17.780 39.510 ;
        RECT 26.030 40.260 26.200 40.430 ;
        RECT 26.950 40.260 27.120 40.430 ;
        RECT 28.580 40.170 28.750 40.340 ;
        RECT 35.870 40.460 36.040 40.630 ;
        RECT 25.520 39.820 25.690 39.990 ;
        RECT 19.560 39.000 19.730 39.170 ;
        RECT 16.510 38.590 16.680 38.760 ;
        RECT 18.150 38.590 18.320 38.760 ;
        RECT 19.060 38.590 19.230 38.760 ;
        RECT 20.670 38.630 20.840 38.800 ;
        RECT 23.360 39.340 23.530 39.510 ;
        RECT 31.780 40.260 31.950 40.430 ;
        RECT 32.700 40.260 32.870 40.430 ;
        RECT 34.330 40.170 34.500 40.340 ;
        RECT 41.620 40.460 41.790 40.630 ;
        RECT 31.270 39.820 31.440 39.990 ;
        RECT 25.310 39.000 25.480 39.170 ;
        RECT 22.260 38.590 22.430 38.760 ;
        RECT 23.900 38.590 24.070 38.760 ;
        RECT 24.810 38.590 24.980 38.760 ;
        RECT 26.420 38.630 26.590 38.800 ;
        RECT 29.110 39.340 29.280 39.510 ;
        RECT 37.530 40.260 37.700 40.430 ;
        RECT 38.450 40.260 38.620 40.430 ;
        RECT 40.080 40.170 40.250 40.340 ;
        RECT 47.370 40.460 47.540 40.630 ;
        RECT 37.020 39.820 37.190 39.990 ;
        RECT 31.060 39.000 31.230 39.170 ;
        RECT 28.010 38.590 28.180 38.760 ;
        RECT 29.650 38.590 29.820 38.760 ;
        RECT 30.560 38.590 30.730 38.760 ;
        RECT 32.170 38.630 32.340 38.800 ;
        RECT 34.860 39.340 35.030 39.510 ;
        RECT 43.280 40.260 43.450 40.430 ;
        RECT 44.200 40.260 44.370 40.430 ;
        RECT 45.830 40.170 46.000 40.340 ;
        RECT 53.120 40.460 53.290 40.630 ;
        RECT 42.770 39.820 42.940 39.990 ;
        RECT 36.810 39.000 36.980 39.170 ;
        RECT 33.760 38.590 33.930 38.760 ;
        RECT 35.400 38.590 35.570 38.760 ;
        RECT 36.310 38.590 36.480 38.760 ;
        RECT 37.920 38.630 38.090 38.800 ;
        RECT 40.610 39.340 40.780 39.510 ;
        RECT 49.030 40.260 49.200 40.430 ;
        RECT 49.950 40.260 50.120 40.430 ;
        RECT 51.580 40.170 51.750 40.340 ;
        RECT 58.870 40.460 59.040 40.630 ;
        RECT 48.520 39.820 48.690 39.990 ;
        RECT 42.560 39.000 42.730 39.170 ;
        RECT 39.510 38.590 39.680 38.760 ;
        RECT 41.150 38.590 41.320 38.760 ;
        RECT 42.060 38.590 42.230 38.760 ;
        RECT 43.670 38.630 43.840 38.800 ;
        RECT 46.360 39.340 46.530 39.510 ;
        RECT 54.780 40.260 54.950 40.430 ;
        RECT 55.700 40.260 55.870 40.430 ;
        RECT 57.330 40.170 57.500 40.340 ;
        RECT 64.620 40.460 64.790 40.630 ;
        RECT 54.270 39.820 54.440 39.990 ;
        RECT 48.310 39.000 48.480 39.170 ;
        RECT 45.260 38.590 45.430 38.760 ;
        RECT 46.900 38.590 47.070 38.760 ;
        RECT 47.810 38.590 47.980 38.760 ;
        RECT 49.420 38.630 49.590 38.800 ;
        RECT 52.110 39.340 52.280 39.510 ;
        RECT 60.530 40.260 60.700 40.430 ;
        RECT 61.450 40.260 61.620 40.430 ;
        RECT 63.080 40.170 63.250 40.340 ;
        RECT 70.370 40.460 70.540 40.630 ;
        RECT 60.020 39.820 60.190 39.990 ;
        RECT 54.060 39.000 54.230 39.170 ;
        RECT 51.010 38.590 51.180 38.760 ;
        RECT 52.650 38.590 52.820 38.760 ;
        RECT 53.560 38.590 53.730 38.760 ;
        RECT 55.170 38.630 55.340 38.800 ;
        RECT 57.860 39.340 58.030 39.510 ;
        RECT 66.280 40.260 66.450 40.430 ;
        RECT 67.200 40.260 67.370 40.430 ;
        RECT 68.830 40.170 69.000 40.340 ;
        RECT 76.120 40.460 76.290 40.630 ;
        RECT 65.770 39.820 65.940 39.990 ;
        RECT 59.810 39.000 59.980 39.170 ;
        RECT 56.760 38.590 56.930 38.760 ;
        RECT 58.400 38.590 58.570 38.760 ;
        RECT 59.310 38.590 59.480 38.760 ;
        RECT 60.920 38.630 61.090 38.800 ;
        RECT 63.610 39.340 63.780 39.510 ;
        RECT 72.030 40.260 72.200 40.430 ;
        RECT 72.950 40.260 73.120 40.430 ;
        RECT 74.580 40.170 74.750 40.340 ;
        RECT 81.870 40.460 82.040 40.630 ;
        RECT 71.520 39.820 71.690 39.990 ;
        RECT 65.560 39.000 65.730 39.170 ;
        RECT 62.510 38.590 62.680 38.760 ;
        RECT 64.150 38.590 64.320 38.760 ;
        RECT 65.060 38.590 65.230 38.760 ;
        RECT 66.670 38.630 66.840 38.800 ;
        RECT 69.360 39.340 69.530 39.510 ;
        RECT 77.780 40.260 77.950 40.430 ;
        RECT 78.700 40.260 78.870 40.430 ;
        RECT 80.330 40.170 80.500 40.340 ;
        RECT 87.620 40.460 87.790 40.630 ;
        RECT 77.270 39.820 77.440 39.990 ;
        RECT 71.310 39.000 71.480 39.170 ;
        RECT 68.260 38.590 68.430 38.760 ;
        RECT 69.900 38.590 70.070 38.760 ;
        RECT 70.810 38.590 70.980 38.760 ;
        RECT 72.420 38.630 72.590 38.800 ;
        RECT 75.110 39.340 75.280 39.510 ;
        RECT 83.530 40.260 83.700 40.430 ;
        RECT 84.450 40.260 84.620 40.430 ;
        RECT 86.080 40.170 86.250 40.340 ;
        RECT 93.370 40.460 93.540 40.630 ;
        RECT 83.020 39.820 83.190 39.990 ;
        RECT 77.060 39.000 77.230 39.170 ;
        RECT 74.010 38.590 74.180 38.760 ;
        RECT 75.650 38.590 75.820 38.760 ;
        RECT 76.560 38.590 76.730 38.760 ;
        RECT 78.170 38.630 78.340 38.800 ;
        RECT 80.860 39.340 81.030 39.510 ;
        RECT 89.280 40.260 89.450 40.430 ;
        RECT 90.200 40.260 90.370 40.430 ;
        RECT 91.830 40.170 92.000 40.340 ;
        RECT 88.770 39.820 88.940 39.990 ;
        RECT 82.810 39.000 82.980 39.170 ;
        RECT 79.760 38.590 79.930 38.760 ;
        RECT 81.400 38.590 81.570 38.760 ;
        RECT 82.310 38.590 82.480 38.760 ;
        RECT 83.920 38.630 84.090 38.800 ;
        RECT 86.610 39.340 86.780 39.510 ;
        RECT 88.560 39.000 88.730 39.170 ;
        RECT 85.510 38.590 85.680 38.760 ;
        RECT 87.150 38.590 87.320 38.760 ;
        RECT 88.060 38.590 88.230 38.760 ;
        RECT 89.670 38.630 89.840 38.800 ;
        RECT 92.360 39.340 92.530 39.510 ;
        RECT 94.310 39.000 94.480 39.170 ;
        RECT 91.260 38.590 91.430 38.760 ;
        RECT 92.900 38.590 93.070 38.760 ;
        RECT 93.810 38.590 93.980 38.760 ;
        RECT 7.120 38.050 7.290 38.220 ;
        RECT 3.030 37.850 3.200 38.020 ;
        RECT 3.950 37.850 4.120 38.020 ;
        RECT 5.580 37.760 5.750 37.930 ;
        RECT 12.870 38.050 13.040 38.220 ;
        RECT 2.520 37.410 2.690 37.580 ;
        RECT 8.780 37.850 8.950 38.020 ;
        RECT 9.700 37.850 9.870 38.020 ;
        RECT 11.330 37.760 11.500 37.930 ;
        RECT 18.620 38.050 18.790 38.220 ;
        RECT 8.270 37.410 8.440 37.580 ;
        RECT 3.420 36.220 3.590 36.390 ;
        RECT 6.110 36.930 6.280 37.100 ;
        RECT 14.530 37.850 14.700 38.020 ;
        RECT 15.450 37.850 15.620 38.020 ;
        RECT 17.080 37.760 17.250 37.930 ;
        RECT 24.370 38.050 24.540 38.220 ;
        RECT 14.020 37.410 14.190 37.580 ;
        RECT 8.060 36.590 8.230 36.760 ;
        RECT 5.010 36.180 5.180 36.350 ;
        RECT 6.650 36.180 6.820 36.350 ;
        RECT 7.560 36.180 7.730 36.350 ;
        RECT 9.170 36.220 9.340 36.390 ;
        RECT 11.860 36.930 12.030 37.100 ;
        RECT 20.280 37.850 20.450 38.020 ;
        RECT 21.200 37.850 21.370 38.020 ;
        RECT 22.830 37.760 23.000 37.930 ;
        RECT 30.120 38.050 30.290 38.220 ;
        RECT 19.770 37.410 19.940 37.580 ;
        RECT 13.810 36.590 13.980 36.760 ;
        RECT 10.760 36.180 10.930 36.350 ;
        RECT 12.400 36.180 12.570 36.350 ;
        RECT 13.310 36.180 13.480 36.350 ;
        RECT 14.920 36.220 15.090 36.390 ;
        RECT 17.610 36.930 17.780 37.100 ;
        RECT 26.030 37.850 26.200 38.020 ;
        RECT 26.950 37.850 27.120 38.020 ;
        RECT 28.580 37.760 28.750 37.930 ;
        RECT 35.870 38.050 36.040 38.220 ;
        RECT 25.520 37.410 25.690 37.580 ;
        RECT 19.560 36.590 19.730 36.760 ;
        RECT 16.510 36.180 16.680 36.350 ;
        RECT 18.150 36.180 18.320 36.350 ;
        RECT 19.060 36.180 19.230 36.350 ;
        RECT 20.670 36.220 20.840 36.390 ;
        RECT 23.360 36.930 23.530 37.100 ;
        RECT 31.780 37.850 31.950 38.020 ;
        RECT 32.700 37.850 32.870 38.020 ;
        RECT 34.330 37.760 34.500 37.930 ;
        RECT 41.620 38.050 41.790 38.220 ;
        RECT 31.270 37.410 31.440 37.580 ;
        RECT 25.310 36.590 25.480 36.760 ;
        RECT 22.260 36.180 22.430 36.350 ;
        RECT 23.900 36.180 24.070 36.350 ;
        RECT 24.810 36.180 24.980 36.350 ;
        RECT 26.420 36.220 26.590 36.390 ;
        RECT 29.110 36.930 29.280 37.100 ;
        RECT 37.530 37.850 37.700 38.020 ;
        RECT 38.450 37.850 38.620 38.020 ;
        RECT 40.080 37.760 40.250 37.930 ;
        RECT 47.370 38.050 47.540 38.220 ;
        RECT 37.020 37.410 37.190 37.580 ;
        RECT 31.060 36.590 31.230 36.760 ;
        RECT 28.010 36.180 28.180 36.350 ;
        RECT 29.650 36.180 29.820 36.350 ;
        RECT 30.560 36.180 30.730 36.350 ;
        RECT 32.170 36.220 32.340 36.390 ;
        RECT 34.860 36.930 35.030 37.100 ;
        RECT 43.280 37.850 43.450 38.020 ;
        RECT 44.200 37.850 44.370 38.020 ;
        RECT 45.830 37.760 46.000 37.930 ;
        RECT 53.120 38.050 53.290 38.220 ;
        RECT 42.770 37.410 42.940 37.580 ;
        RECT 36.810 36.590 36.980 36.760 ;
        RECT 33.760 36.180 33.930 36.350 ;
        RECT 35.400 36.180 35.570 36.350 ;
        RECT 36.310 36.180 36.480 36.350 ;
        RECT 37.920 36.220 38.090 36.390 ;
        RECT 40.610 36.930 40.780 37.100 ;
        RECT 49.030 37.850 49.200 38.020 ;
        RECT 49.950 37.850 50.120 38.020 ;
        RECT 51.580 37.760 51.750 37.930 ;
        RECT 58.870 38.050 59.040 38.220 ;
        RECT 48.520 37.410 48.690 37.580 ;
        RECT 42.560 36.590 42.730 36.760 ;
        RECT 39.510 36.180 39.680 36.350 ;
        RECT 41.150 36.180 41.320 36.350 ;
        RECT 42.060 36.180 42.230 36.350 ;
        RECT 43.670 36.220 43.840 36.390 ;
        RECT 46.360 36.930 46.530 37.100 ;
        RECT 54.780 37.850 54.950 38.020 ;
        RECT 55.700 37.850 55.870 38.020 ;
        RECT 57.330 37.760 57.500 37.930 ;
        RECT 64.620 38.050 64.790 38.220 ;
        RECT 54.270 37.410 54.440 37.580 ;
        RECT 48.310 36.590 48.480 36.760 ;
        RECT 45.260 36.180 45.430 36.350 ;
        RECT 46.900 36.180 47.070 36.350 ;
        RECT 47.810 36.180 47.980 36.350 ;
        RECT 49.420 36.220 49.590 36.390 ;
        RECT 52.110 36.930 52.280 37.100 ;
        RECT 60.530 37.850 60.700 38.020 ;
        RECT 61.450 37.850 61.620 38.020 ;
        RECT 63.080 37.760 63.250 37.930 ;
        RECT 70.370 38.050 70.540 38.220 ;
        RECT 60.020 37.410 60.190 37.580 ;
        RECT 54.060 36.590 54.230 36.760 ;
        RECT 51.010 36.180 51.180 36.350 ;
        RECT 52.650 36.180 52.820 36.350 ;
        RECT 53.560 36.180 53.730 36.350 ;
        RECT 55.170 36.220 55.340 36.390 ;
        RECT 57.860 36.930 58.030 37.100 ;
        RECT 66.280 37.850 66.450 38.020 ;
        RECT 67.200 37.850 67.370 38.020 ;
        RECT 68.830 37.760 69.000 37.930 ;
        RECT 76.120 38.050 76.290 38.220 ;
        RECT 65.770 37.410 65.940 37.580 ;
        RECT 59.810 36.590 59.980 36.760 ;
        RECT 56.760 36.180 56.930 36.350 ;
        RECT 58.400 36.180 58.570 36.350 ;
        RECT 59.310 36.180 59.480 36.350 ;
        RECT 60.920 36.220 61.090 36.390 ;
        RECT 63.610 36.930 63.780 37.100 ;
        RECT 72.030 37.850 72.200 38.020 ;
        RECT 72.950 37.850 73.120 38.020 ;
        RECT 74.580 37.760 74.750 37.930 ;
        RECT 81.870 38.050 82.040 38.220 ;
        RECT 71.520 37.410 71.690 37.580 ;
        RECT 65.560 36.590 65.730 36.760 ;
        RECT 62.510 36.180 62.680 36.350 ;
        RECT 64.150 36.180 64.320 36.350 ;
        RECT 65.060 36.180 65.230 36.350 ;
        RECT 66.670 36.220 66.840 36.390 ;
        RECT 69.360 36.930 69.530 37.100 ;
        RECT 77.780 37.850 77.950 38.020 ;
        RECT 78.700 37.850 78.870 38.020 ;
        RECT 80.330 37.760 80.500 37.930 ;
        RECT 87.620 38.050 87.790 38.220 ;
        RECT 77.270 37.410 77.440 37.580 ;
        RECT 71.310 36.590 71.480 36.760 ;
        RECT 68.260 36.180 68.430 36.350 ;
        RECT 69.900 36.180 70.070 36.350 ;
        RECT 70.810 36.180 70.980 36.350 ;
        RECT 72.420 36.220 72.590 36.390 ;
        RECT 75.110 36.930 75.280 37.100 ;
        RECT 83.530 37.850 83.700 38.020 ;
        RECT 84.450 37.850 84.620 38.020 ;
        RECT 86.080 37.760 86.250 37.930 ;
        RECT 93.370 38.050 93.540 38.220 ;
        RECT 83.020 37.410 83.190 37.580 ;
        RECT 77.060 36.590 77.230 36.760 ;
        RECT 74.010 36.180 74.180 36.350 ;
        RECT 75.650 36.180 75.820 36.350 ;
        RECT 76.560 36.180 76.730 36.350 ;
        RECT 78.170 36.220 78.340 36.390 ;
        RECT 80.860 36.930 81.030 37.100 ;
        RECT 89.280 37.850 89.450 38.020 ;
        RECT 90.200 37.850 90.370 38.020 ;
        RECT 91.830 37.760 92.000 37.930 ;
        RECT 88.770 37.410 88.940 37.580 ;
        RECT 82.810 36.590 82.980 36.760 ;
        RECT 79.760 36.180 79.930 36.350 ;
        RECT 81.400 36.180 81.570 36.350 ;
        RECT 82.310 36.180 82.480 36.350 ;
        RECT 83.920 36.220 84.090 36.390 ;
        RECT 86.610 36.930 86.780 37.100 ;
        RECT 88.560 36.590 88.730 36.760 ;
        RECT 85.510 36.180 85.680 36.350 ;
        RECT 87.150 36.180 87.320 36.350 ;
        RECT 88.060 36.180 88.230 36.350 ;
        RECT 89.670 36.220 89.840 36.390 ;
        RECT 92.360 36.930 92.530 37.100 ;
        RECT 94.310 36.590 94.480 36.760 ;
        RECT 91.260 36.180 91.430 36.350 ;
        RECT 92.900 36.180 93.070 36.350 ;
        RECT 93.810 36.180 93.980 36.350 ;
        RECT 7.120 35.640 7.290 35.810 ;
        RECT 3.030 35.440 3.200 35.610 ;
        RECT 3.950 35.440 4.120 35.610 ;
        RECT 5.580 35.350 5.750 35.520 ;
        RECT 12.870 35.640 13.040 35.810 ;
        RECT 2.520 35.000 2.690 35.170 ;
        RECT 8.780 35.440 8.950 35.610 ;
        RECT 9.700 35.440 9.870 35.610 ;
        RECT 11.330 35.350 11.500 35.520 ;
        RECT 18.620 35.640 18.790 35.810 ;
        RECT 8.270 35.000 8.440 35.170 ;
        RECT 3.420 33.810 3.590 33.980 ;
        RECT 6.110 34.520 6.280 34.690 ;
        RECT 14.530 35.440 14.700 35.610 ;
        RECT 15.450 35.440 15.620 35.610 ;
        RECT 17.080 35.350 17.250 35.520 ;
        RECT 24.370 35.640 24.540 35.810 ;
        RECT 14.020 35.000 14.190 35.170 ;
        RECT 8.060 34.180 8.230 34.350 ;
        RECT 5.010 33.770 5.180 33.940 ;
        RECT 6.650 33.770 6.820 33.940 ;
        RECT 7.560 33.770 7.730 33.940 ;
        RECT 9.170 33.810 9.340 33.980 ;
        RECT 11.860 34.520 12.030 34.690 ;
        RECT 20.280 35.440 20.450 35.610 ;
        RECT 21.200 35.440 21.370 35.610 ;
        RECT 22.830 35.350 23.000 35.520 ;
        RECT 30.120 35.640 30.290 35.810 ;
        RECT 19.770 35.000 19.940 35.170 ;
        RECT 13.810 34.180 13.980 34.350 ;
        RECT 10.760 33.770 10.930 33.940 ;
        RECT 12.400 33.770 12.570 33.940 ;
        RECT 13.310 33.770 13.480 33.940 ;
        RECT 14.920 33.810 15.090 33.980 ;
        RECT 17.610 34.520 17.780 34.690 ;
        RECT 26.030 35.440 26.200 35.610 ;
        RECT 26.950 35.440 27.120 35.610 ;
        RECT 28.580 35.350 28.750 35.520 ;
        RECT 35.870 35.640 36.040 35.810 ;
        RECT 25.520 35.000 25.690 35.170 ;
        RECT 19.560 34.180 19.730 34.350 ;
        RECT 16.510 33.770 16.680 33.940 ;
        RECT 18.150 33.770 18.320 33.940 ;
        RECT 19.060 33.770 19.230 33.940 ;
        RECT 20.670 33.810 20.840 33.980 ;
        RECT 23.360 34.520 23.530 34.690 ;
        RECT 31.780 35.440 31.950 35.610 ;
        RECT 32.700 35.440 32.870 35.610 ;
        RECT 34.330 35.350 34.500 35.520 ;
        RECT 41.620 35.640 41.790 35.810 ;
        RECT 31.270 35.000 31.440 35.170 ;
        RECT 25.310 34.180 25.480 34.350 ;
        RECT 22.260 33.770 22.430 33.940 ;
        RECT 23.900 33.770 24.070 33.940 ;
        RECT 24.810 33.770 24.980 33.940 ;
        RECT 26.420 33.810 26.590 33.980 ;
        RECT 29.110 34.520 29.280 34.690 ;
        RECT 37.530 35.440 37.700 35.610 ;
        RECT 38.450 35.440 38.620 35.610 ;
        RECT 40.080 35.350 40.250 35.520 ;
        RECT 47.370 35.640 47.540 35.810 ;
        RECT 37.020 35.000 37.190 35.170 ;
        RECT 31.060 34.180 31.230 34.350 ;
        RECT 28.010 33.770 28.180 33.940 ;
        RECT 29.650 33.770 29.820 33.940 ;
        RECT 30.560 33.770 30.730 33.940 ;
        RECT 32.170 33.810 32.340 33.980 ;
        RECT 34.860 34.520 35.030 34.690 ;
        RECT 43.280 35.440 43.450 35.610 ;
        RECT 44.200 35.440 44.370 35.610 ;
        RECT 45.830 35.350 46.000 35.520 ;
        RECT 53.120 35.640 53.290 35.810 ;
        RECT 42.770 35.000 42.940 35.170 ;
        RECT 36.810 34.180 36.980 34.350 ;
        RECT 33.760 33.770 33.930 33.940 ;
        RECT 35.400 33.770 35.570 33.940 ;
        RECT 36.310 33.770 36.480 33.940 ;
        RECT 37.920 33.810 38.090 33.980 ;
        RECT 40.610 34.520 40.780 34.690 ;
        RECT 49.030 35.440 49.200 35.610 ;
        RECT 49.950 35.440 50.120 35.610 ;
        RECT 51.580 35.350 51.750 35.520 ;
        RECT 58.870 35.640 59.040 35.810 ;
        RECT 48.520 35.000 48.690 35.170 ;
        RECT 42.560 34.180 42.730 34.350 ;
        RECT 39.510 33.770 39.680 33.940 ;
        RECT 41.150 33.770 41.320 33.940 ;
        RECT 42.060 33.770 42.230 33.940 ;
        RECT 43.670 33.810 43.840 33.980 ;
        RECT 46.360 34.520 46.530 34.690 ;
        RECT 54.780 35.440 54.950 35.610 ;
        RECT 55.700 35.440 55.870 35.610 ;
        RECT 57.330 35.350 57.500 35.520 ;
        RECT 64.620 35.640 64.790 35.810 ;
        RECT 54.270 35.000 54.440 35.170 ;
        RECT 48.310 34.180 48.480 34.350 ;
        RECT 45.260 33.770 45.430 33.940 ;
        RECT 46.900 33.770 47.070 33.940 ;
        RECT 47.810 33.770 47.980 33.940 ;
        RECT 49.420 33.810 49.590 33.980 ;
        RECT 52.110 34.520 52.280 34.690 ;
        RECT 60.530 35.440 60.700 35.610 ;
        RECT 61.450 35.440 61.620 35.610 ;
        RECT 63.080 35.350 63.250 35.520 ;
        RECT 70.370 35.640 70.540 35.810 ;
        RECT 60.020 35.000 60.190 35.170 ;
        RECT 54.060 34.180 54.230 34.350 ;
        RECT 51.010 33.770 51.180 33.940 ;
        RECT 52.650 33.770 52.820 33.940 ;
        RECT 53.560 33.770 53.730 33.940 ;
        RECT 55.170 33.810 55.340 33.980 ;
        RECT 57.860 34.520 58.030 34.690 ;
        RECT 66.280 35.440 66.450 35.610 ;
        RECT 67.200 35.440 67.370 35.610 ;
        RECT 68.830 35.350 69.000 35.520 ;
        RECT 76.120 35.640 76.290 35.810 ;
        RECT 65.770 35.000 65.940 35.170 ;
        RECT 59.810 34.180 59.980 34.350 ;
        RECT 56.760 33.770 56.930 33.940 ;
        RECT 58.400 33.770 58.570 33.940 ;
        RECT 59.310 33.770 59.480 33.940 ;
        RECT 60.920 33.810 61.090 33.980 ;
        RECT 63.610 34.520 63.780 34.690 ;
        RECT 72.030 35.440 72.200 35.610 ;
        RECT 72.950 35.440 73.120 35.610 ;
        RECT 74.580 35.350 74.750 35.520 ;
        RECT 81.870 35.640 82.040 35.810 ;
        RECT 71.520 35.000 71.690 35.170 ;
        RECT 65.560 34.180 65.730 34.350 ;
        RECT 62.510 33.770 62.680 33.940 ;
        RECT 64.150 33.770 64.320 33.940 ;
        RECT 65.060 33.770 65.230 33.940 ;
        RECT 66.670 33.810 66.840 33.980 ;
        RECT 69.360 34.520 69.530 34.690 ;
        RECT 77.780 35.440 77.950 35.610 ;
        RECT 78.700 35.440 78.870 35.610 ;
        RECT 80.330 35.350 80.500 35.520 ;
        RECT 87.620 35.640 87.790 35.810 ;
        RECT 77.270 35.000 77.440 35.170 ;
        RECT 71.310 34.180 71.480 34.350 ;
        RECT 68.260 33.770 68.430 33.940 ;
        RECT 69.900 33.770 70.070 33.940 ;
        RECT 70.810 33.770 70.980 33.940 ;
        RECT 72.420 33.810 72.590 33.980 ;
        RECT 75.110 34.520 75.280 34.690 ;
        RECT 83.530 35.440 83.700 35.610 ;
        RECT 84.450 35.440 84.620 35.610 ;
        RECT 86.080 35.350 86.250 35.520 ;
        RECT 93.370 35.640 93.540 35.810 ;
        RECT 83.020 35.000 83.190 35.170 ;
        RECT 77.060 34.180 77.230 34.350 ;
        RECT 74.010 33.770 74.180 33.940 ;
        RECT 75.650 33.770 75.820 33.940 ;
        RECT 76.560 33.770 76.730 33.940 ;
        RECT 78.170 33.810 78.340 33.980 ;
        RECT 80.860 34.520 81.030 34.690 ;
        RECT 89.280 35.440 89.450 35.610 ;
        RECT 90.200 35.440 90.370 35.610 ;
        RECT 91.830 35.350 92.000 35.520 ;
        RECT 88.770 35.000 88.940 35.170 ;
        RECT 82.810 34.180 82.980 34.350 ;
        RECT 79.760 33.770 79.930 33.940 ;
        RECT 81.400 33.770 81.570 33.940 ;
        RECT 82.310 33.770 82.480 33.940 ;
        RECT 83.920 33.810 84.090 33.980 ;
        RECT 86.610 34.520 86.780 34.690 ;
        RECT 88.560 34.180 88.730 34.350 ;
        RECT 85.510 33.770 85.680 33.940 ;
        RECT 87.150 33.770 87.320 33.940 ;
        RECT 88.060 33.770 88.230 33.940 ;
        RECT 89.670 33.810 89.840 33.980 ;
        RECT 92.360 34.520 92.530 34.690 ;
        RECT 94.310 34.180 94.480 34.350 ;
        RECT 91.260 33.770 91.430 33.940 ;
        RECT 92.900 33.770 93.070 33.940 ;
        RECT 93.810 33.770 93.980 33.940 ;
        RECT 7.120 33.230 7.290 33.400 ;
        RECT 3.030 33.030 3.200 33.200 ;
        RECT 3.950 33.030 4.120 33.200 ;
        RECT 5.580 32.940 5.750 33.110 ;
        RECT 12.870 33.230 13.040 33.400 ;
        RECT 2.520 32.590 2.690 32.760 ;
        RECT 8.780 33.030 8.950 33.200 ;
        RECT 9.700 33.030 9.870 33.200 ;
        RECT 11.330 32.940 11.500 33.110 ;
        RECT 18.620 33.230 18.790 33.400 ;
        RECT 8.270 32.590 8.440 32.760 ;
        RECT 3.420 31.400 3.590 31.570 ;
        RECT 6.110 32.110 6.280 32.280 ;
        RECT 14.530 33.030 14.700 33.200 ;
        RECT 15.450 33.030 15.620 33.200 ;
        RECT 17.080 32.940 17.250 33.110 ;
        RECT 24.370 33.230 24.540 33.400 ;
        RECT 14.020 32.590 14.190 32.760 ;
        RECT 8.060 31.770 8.230 31.940 ;
        RECT 5.010 31.360 5.180 31.530 ;
        RECT 6.650 31.360 6.820 31.530 ;
        RECT 7.560 31.360 7.730 31.530 ;
        RECT 9.170 31.400 9.340 31.570 ;
        RECT 11.860 32.110 12.030 32.280 ;
        RECT 20.280 33.030 20.450 33.200 ;
        RECT 21.200 33.030 21.370 33.200 ;
        RECT 22.830 32.940 23.000 33.110 ;
        RECT 30.120 33.230 30.290 33.400 ;
        RECT 19.770 32.590 19.940 32.760 ;
        RECT 13.810 31.770 13.980 31.940 ;
        RECT 10.760 31.360 10.930 31.530 ;
        RECT 12.400 31.360 12.570 31.530 ;
        RECT 13.310 31.360 13.480 31.530 ;
        RECT 14.920 31.400 15.090 31.570 ;
        RECT 17.610 32.110 17.780 32.280 ;
        RECT 26.030 33.030 26.200 33.200 ;
        RECT 26.950 33.030 27.120 33.200 ;
        RECT 28.580 32.940 28.750 33.110 ;
        RECT 35.870 33.230 36.040 33.400 ;
        RECT 25.520 32.590 25.690 32.760 ;
        RECT 19.560 31.770 19.730 31.940 ;
        RECT 16.510 31.360 16.680 31.530 ;
        RECT 18.150 31.360 18.320 31.530 ;
        RECT 19.060 31.360 19.230 31.530 ;
        RECT 20.670 31.400 20.840 31.570 ;
        RECT 23.360 32.110 23.530 32.280 ;
        RECT 31.780 33.030 31.950 33.200 ;
        RECT 32.700 33.030 32.870 33.200 ;
        RECT 34.330 32.940 34.500 33.110 ;
        RECT 41.620 33.230 41.790 33.400 ;
        RECT 31.270 32.590 31.440 32.760 ;
        RECT 25.310 31.770 25.480 31.940 ;
        RECT 22.260 31.360 22.430 31.530 ;
        RECT 23.900 31.360 24.070 31.530 ;
        RECT 24.810 31.360 24.980 31.530 ;
        RECT 26.420 31.400 26.590 31.570 ;
        RECT 29.110 32.110 29.280 32.280 ;
        RECT 37.530 33.030 37.700 33.200 ;
        RECT 38.450 33.030 38.620 33.200 ;
        RECT 40.080 32.940 40.250 33.110 ;
        RECT 47.370 33.230 47.540 33.400 ;
        RECT 37.020 32.590 37.190 32.760 ;
        RECT 31.060 31.770 31.230 31.940 ;
        RECT 28.010 31.360 28.180 31.530 ;
        RECT 29.650 31.360 29.820 31.530 ;
        RECT 30.560 31.360 30.730 31.530 ;
        RECT 32.170 31.400 32.340 31.570 ;
        RECT 34.860 32.110 35.030 32.280 ;
        RECT 43.280 33.030 43.450 33.200 ;
        RECT 44.200 33.030 44.370 33.200 ;
        RECT 45.830 32.940 46.000 33.110 ;
        RECT 53.120 33.230 53.290 33.400 ;
        RECT 42.770 32.590 42.940 32.760 ;
        RECT 36.810 31.770 36.980 31.940 ;
        RECT 33.760 31.360 33.930 31.530 ;
        RECT 35.400 31.360 35.570 31.530 ;
        RECT 36.310 31.360 36.480 31.530 ;
        RECT 37.920 31.400 38.090 31.570 ;
        RECT 40.610 32.110 40.780 32.280 ;
        RECT 49.030 33.030 49.200 33.200 ;
        RECT 49.950 33.030 50.120 33.200 ;
        RECT 51.580 32.940 51.750 33.110 ;
        RECT 58.870 33.230 59.040 33.400 ;
        RECT 48.520 32.590 48.690 32.760 ;
        RECT 42.560 31.770 42.730 31.940 ;
        RECT 39.510 31.360 39.680 31.530 ;
        RECT 41.150 31.360 41.320 31.530 ;
        RECT 42.060 31.360 42.230 31.530 ;
        RECT 43.670 31.400 43.840 31.570 ;
        RECT 46.360 32.110 46.530 32.280 ;
        RECT 54.780 33.030 54.950 33.200 ;
        RECT 55.700 33.030 55.870 33.200 ;
        RECT 57.330 32.940 57.500 33.110 ;
        RECT 64.620 33.230 64.790 33.400 ;
        RECT 54.270 32.590 54.440 32.760 ;
        RECT 48.310 31.770 48.480 31.940 ;
        RECT 45.260 31.360 45.430 31.530 ;
        RECT 46.900 31.360 47.070 31.530 ;
        RECT 47.810 31.360 47.980 31.530 ;
        RECT 49.420 31.400 49.590 31.570 ;
        RECT 52.110 32.110 52.280 32.280 ;
        RECT 60.530 33.030 60.700 33.200 ;
        RECT 61.450 33.030 61.620 33.200 ;
        RECT 63.080 32.940 63.250 33.110 ;
        RECT 70.370 33.230 70.540 33.400 ;
        RECT 60.020 32.590 60.190 32.760 ;
        RECT 54.060 31.770 54.230 31.940 ;
        RECT 51.010 31.360 51.180 31.530 ;
        RECT 52.650 31.360 52.820 31.530 ;
        RECT 53.560 31.360 53.730 31.530 ;
        RECT 55.170 31.400 55.340 31.570 ;
        RECT 57.860 32.110 58.030 32.280 ;
        RECT 66.280 33.030 66.450 33.200 ;
        RECT 67.200 33.030 67.370 33.200 ;
        RECT 68.830 32.940 69.000 33.110 ;
        RECT 76.120 33.230 76.290 33.400 ;
        RECT 65.770 32.590 65.940 32.760 ;
        RECT 59.810 31.770 59.980 31.940 ;
        RECT 56.760 31.360 56.930 31.530 ;
        RECT 58.400 31.360 58.570 31.530 ;
        RECT 59.310 31.360 59.480 31.530 ;
        RECT 60.920 31.400 61.090 31.570 ;
        RECT 63.610 32.110 63.780 32.280 ;
        RECT 72.030 33.030 72.200 33.200 ;
        RECT 72.950 33.030 73.120 33.200 ;
        RECT 74.580 32.940 74.750 33.110 ;
        RECT 81.870 33.230 82.040 33.400 ;
        RECT 71.520 32.590 71.690 32.760 ;
        RECT 65.560 31.770 65.730 31.940 ;
        RECT 62.510 31.360 62.680 31.530 ;
        RECT 64.150 31.360 64.320 31.530 ;
        RECT 65.060 31.360 65.230 31.530 ;
        RECT 66.670 31.400 66.840 31.570 ;
        RECT 69.360 32.110 69.530 32.280 ;
        RECT 77.780 33.030 77.950 33.200 ;
        RECT 78.700 33.030 78.870 33.200 ;
        RECT 80.330 32.940 80.500 33.110 ;
        RECT 87.620 33.230 87.790 33.400 ;
        RECT 77.270 32.590 77.440 32.760 ;
        RECT 71.310 31.770 71.480 31.940 ;
        RECT 68.260 31.360 68.430 31.530 ;
        RECT 69.900 31.360 70.070 31.530 ;
        RECT 70.810 31.360 70.980 31.530 ;
        RECT 72.420 31.400 72.590 31.570 ;
        RECT 75.110 32.110 75.280 32.280 ;
        RECT 83.530 33.030 83.700 33.200 ;
        RECT 84.450 33.030 84.620 33.200 ;
        RECT 86.080 32.940 86.250 33.110 ;
        RECT 93.370 33.230 93.540 33.400 ;
        RECT 83.020 32.590 83.190 32.760 ;
        RECT 77.060 31.770 77.230 31.940 ;
        RECT 74.010 31.360 74.180 31.530 ;
        RECT 75.650 31.360 75.820 31.530 ;
        RECT 76.560 31.360 76.730 31.530 ;
        RECT 78.170 31.400 78.340 31.570 ;
        RECT 80.860 32.110 81.030 32.280 ;
        RECT 89.280 33.030 89.450 33.200 ;
        RECT 90.200 33.030 90.370 33.200 ;
        RECT 91.830 32.940 92.000 33.110 ;
        RECT 88.770 32.590 88.940 32.760 ;
        RECT 82.810 31.770 82.980 31.940 ;
        RECT 79.760 31.360 79.930 31.530 ;
        RECT 81.400 31.360 81.570 31.530 ;
        RECT 82.310 31.360 82.480 31.530 ;
        RECT 83.920 31.400 84.090 31.570 ;
        RECT 86.610 32.110 86.780 32.280 ;
        RECT 88.560 31.770 88.730 31.940 ;
        RECT 85.510 31.360 85.680 31.530 ;
        RECT 87.150 31.360 87.320 31.530 ;
        RECT 88.060 31.360 88.230 31.530 ;
        RECT 89.670 31.400 89.840 31.570 ;
        RECT 92.360 32.110 92.530 32.280 ;
        RECT 94.310 31.770 94.480 31.940 ;
        RECT 91.260 31.360 91.430 31.530 ;
        RECT 92.900 31.360 93.070 31.530 ;
        RECT 93.810 31.360 93.980 31.530 ;
        RECT 7.120 30.820 7.290 30.990 ;
        RECT 3.030 30.620 3.200 30.790 ;
        RECT 3.950 30.620 4.120 30.790 ;
        RECT 5.580 30.530 5.750 30.700 ;
        RECT 12.870 30.820 13.040 30.990 ;
        RECT 2.520 30.180 2.690 30.350 ;
        RECT 8.780 30.620 8.950 30.790 ;
        RECT 9.700 30.620 9.870 30.790 ;
        RECT 11.330 30.530 11.500 30.700 ;
        RECT 18.620 30.820 18.790 30.990 ;
        RECT 8.270 30.180 8.440 30.350 ;
        RECT 3.420 28.990 3.590 29.160 ;
        RECT 6.110 29.700 6.280 29.870 ;
        RECT 14.530 30.620 14.700 30.790 ;
        RECT 15.450 30.620 15.620 30.790 ;
        RECT 17.080 30.530 17.250 30.700 ;
        RECT 24.370 30.820 24.540 30.990 ;
        RECT 14.020 30.180 14.190 30.350 ;
        RECT 8.060 29.360 8.230 29.530 ;
        RECT 5.010 28.950 5.180 29.120 ;
        RECT 6.650 28.950 6.820 29.120 ;
        RECT 7.560 28.950 7.730 29.120 ;
        RECT 7.120 28.090 7.290 28.260 ;
        RECT 9.170 28.990 9.340 29.160 ;
        RECT 11.860 29.700 12.030 29.870 ;
        RECT 20.280 30.620 20.450 30.790 ;
        RECT 21.200 30.620 21.370 30.790 ;
        RECT 22.830 30.530 23.000 30.700 ;
        RECT 30.120 30.820 30.290 30.990 ;
        RECT 19.770 30.180 19.940 30.350 ;
        RECT 13.810 29.360 13.980 29.530 ;
        RECT 10.760 28.950 10.930 29.120 ;
        RECT 12.400 28.950 12.570 29.120 ;
        RECT 13.310 28.950 13.480 29.120 ;
        RECT 3.030 27.810 3.200 27.980 ;
        RECT 3.950 27.810 4.120 27.980 ;
        RECT 5.580 27.720 5.750 27.890 ;
        RECT 12.870 28.090 13.040 28.260 ;
        RECT 14.920 28.990 15.090 29.160 ;
        RECT 17.610 29.700 17.780 29.870 ;
        RECT 26.030 30.620 26.200 30.790 ;
        RECT 26.950 30.620 27.120 30.790 ;
        RECT 28.580 30.530 28.750 30.700 ;
        RECT 35.870 30.820 36.040 30.990 ;
        RECT 25.520 30.180 25.690 30.350 ;
        RECT 19.560 29.360 19.730 29.530 ;
        RECT 16.510 28.950 16.680 29.120 ;
        RECT 18.150 28.950 18.320 29.120 ;
        RECT 19.060 28.950 19.230 29.120 ;
        RECT 2.520 27.370 2.690 27.540 ;
        RECT 8.780 27.810 8.950 27.980 ;
        RECT 9.700 27.810 9.870 27.980 ;
        RECT 11.330 27.720 11.500 27.890 ;
        RECT 18.620 28.090 18.790 28.260 ;
        RECT 20.670 28.990 20.840 29.160 ;
        RECT 23.360 29.700 23.530 29.870 ;
        RECT 31.780 30.620 31.950 30.790 ;
        RECT 32.700 30.620 32.870 30.790 ;
        RECT 34.330 30.530 34.500 30.700 ;
        RECT 41.620 30.820 41.790 30.990 ;
        RECT 31.270 30.180 31.440 30.350 ;
        RECT 25.310 29.360 25.480 29.530 ;
        RECT 22.260 28.950 22.430 29.120 ;
        RECT 23.900 28.950 24.070 29.120 ;
        RECT 24.810 28.950 24.980 29.120 ;
        RECT 8.270 27.370 8.440 27.540 ;
        RECT 3.420 26.180 3.590 26.350 ;
        RECT 6.110 26.890 6.280 27.060 ;
        RECT 14.530 27.810 14.700 27.980 ;
        RECT 15.450 27.810 15.620 27.980 ;
        RECT 17.080 27.720 17.250 27.890 ;
        RECT 24.370 28.090 24.540 28.260 ;
        RECT 26.420 28.990 26.590 29.160 ;
        RECT 29.110 29.700 29.280 29.870 ;
        RECT 37.530 30.620 37.700 30.790 ;
        RECT 38.450 30.620 38.620 30.790 ;
        RECT 40.080 30.530 40.250 30.700 ;
        RECT 47.370 30.820 47.540 30.990 ;
        RECT 37.020 30.180 37.190 30.350 ;
        RECT 31.060 29.360 31.230 29.530 ;
        RECT 28.010 28.950 28.180 29.120 ;
        RECT 29.650 28.950 29.820 29.120 ;
        RECT 30.560 28.950 30.730 29.120 ;
        RECT 14.020 27.370 14.190 27.540 ;
        RECT 8.060 26.550 8.230 26.720 ;
        RECT 5.010 26.140 5.180 26.310 ;
        RECT 6.650 26.140 6.820 26.310 ;
        RECT 7.560 26.140 7.730 26.310 ;
        RECT 9.170 26.180 9.340 26.350 ;
        RECT 11.860 26.890 12.030 27.060 ;
        RECT 20.280 27.810 20.450 27.980 ;
        RECT 21.200 27.810 21.370 27.980 ;
        RECT 22.830 27.720 23.000 27.890 ;
        RECT 30.120 28.090 30.290 28.260 ;
        RECT 32.170 28.990 32.340 29.160 ;
        RECT 34.860 29.700 35.030 29.870 ;
        RECT 43.280 30.620 43.450 30.790 ;
        RECT 44.200 30.620 44.370 30.790 ;
        RECT 45.830 30.530 46.000 30.700 ;
        RECT 53.120 30.820 53.290 30.990 ;
        RECT 42.770 30.180 42.940 30.350 ;
        RECT 36.810 29.360 36.980 29.530 ;
        RECT 33.760 28.950 33.930 29.120 ;
        RECT 35.400 28.950 35.570 29.120 ;
        RECT 36.310 28.950 36.480 29.120 ;
        RECT 19.770 27.370 19.940 27.540 ;
        RECT 13.810 26.550 13.980 26.720 ;
        RECT 10.760 26.140 10.930 26.310 ;
        RECT 12.400 26.140 12.570 26.310 ;
        RECT 13.310 26.140 13.480 26.310 ;
        RECT 14.920 26.180 15.090 26.350 ;
        RECT 17.610 26.890 17.780 27.060 ;
        RECT 26.030 27.810 26.200 27.980 ;
        RECT 26.950 27.810 27.120 27.980 ;
        RECT 28.580 27.720 28.750 27.890 ;
        RECT 35.870 28.090 36.040 28.260 ;
        RECT 37.920 28.990 38.090 29.160 ;
        RECT 40.610 29.700 40.780 29.870 ;
        RECT 49.030 30.620 49.200 30.790 ;
        RECT 49.950 30.620 50.120 30.790 ;
        RECT 51.580 30.530 51.750 30.700 ;
        RECT 58.870 30.820 59.040 30.990 ;
        RECT 48.520 30.180 48.690 30.350 ;
        RECT 42.560 29.360 42.730 29.530 ;
        RECT 39.510 28.950 39.680 29.120 ;
        RECT 41.150 28.950 41.320 29.120 ;
        RECT 42.060 28.950 42.230 29.120 ;
        RECT 25.520 27.370 25.690 27.540 ;
        RECT 19.560 26.550 19.730 26.720 ;
        RECT 16.510 26.140 16.680 26.310 ;
        RECT 18.150 26.140 18.320 26.310 ;
        RECT 19.060 26.140 19.230 26.310 ;
        RECT 20.670 26.180 20.840 26.350 ;
        RECT 23.360 26.890 23.530 27.060 ;
        RECT 31.780 27.810 31.950 27.980 ;
        RECT 32.700 27.810 32.870 27.980 ;
        RECT 34.330 27.720 34.500 27.890 ;
        RECT 41.620 28.090 41.790 28.260 ;
        RECT 43.670 28.990 43.840 29.160 ;
        RECT 46.360 29.700 46.530 29.870 ;
        RECT 54.780 30.620 54.950 30.790 ;
        RECT 55.700 30.620 55.870 30.790 ;
        RECT 57.330 30.530 57.500 30.700 ;
        RECT 64.620 30.820 64.790 30.990 ;
        RECT 54.270 30.180 54.440 30.350 ;
        RECT 48.310 29.360 48.480 29.530 ;
        RECT 45.260 28.950 45.430 29.120 ;
        RECT 46.900 28.950 47.070 29.120 ;
        RECT 47.810 28.950 47.980 29.120 ;
        RECT 31.270 27.370 31.440 27.540 ;
        RECT 25.310 26.550 25.480 26.720 ;
        RECT 22.260 26.140 22.430 26.310 ;
        RECT 23.900 26.140 24.070 26.310 ;
        RECT 24.810 26.140 24.980 26.310 ;
        RECT 26.420 26.180 26.590 26.350 ;
        RECT 29.110 26.890 29.280 27.060 ;
        RECT 37.530 27.810 37.700 27.980 ;
        RECT 38.450 27.810 38.620 27.980 ;
        RECT 40.080 27.720 40.250 27.890 ;
        RECT 47.370 28.090 47.540 28.260 ;
        RECT 49.420 28.990 49.590 29.160 ;
        RECT 52.110 29.700 52.280 29.870 ;
        RECT 60.530 30.620 60.700 30.790 ;
        RECT 61.450 30.620 61.620 30.790 ;
        RECT 63.080 30.530 63.250 30.700 ;
        RECT 70.370 30.820 70.540 30.990 ;
        RECT 60.020 30.180 60.190 30.350 ;
        RECT 54.060 29.360 54.230 29.530 ;
        RECT 51.010 28.950 51.180 29.120 ;
        RECT 52.650 28.950 52.820 29.120 ;
        RECT 53.560 28.950 53.730 29.120 ;
        RECT 37.020 27.370 37.190 27.540 ;
        RECT 31.060 26.550 31.230 26.720 ;
        RECT 28.010 26.140 28.180 26.310 ;
        RECT 29.650 26.140 29.820 26.310 ;
        RECT 30.560 26.140 30.730 26.310 ;
        RECT 32.170 26.180 32.340 26.350 ;
        RECT 34.860 26.890 35.030 27.060 ;
        RECT 43.280 27.810 43.450 27.980 ;
        RECT 44.200 27.810 44.370 27.980 ;
        RECT 45.830 27.720 46.000 27.890 ;
        RECT 53.120 28.090 53.290 28.260 ;
        RECT 55.170 28.990 55.340 29.160 ;
        RECT 57.860 29.700 58.030 29.870 ;
        RECT 66.280 30.620 66.450 30.790 ;
        RECT 67.200 30.620 67.370 30.790 ;
        RECT 68.830 30.530 69.000 30.700 ;
        RECT 76.120 30.820 76.290 30.990 ;
        RECT 65.770 30.180 65.940 30.350 ;
        RECT 59.810 29.360 59.980 29.530 ;
        RECT 56.760 28.950 56.930 29.120 ;
        RECT 58.400 28.950 58.570 29.120 ;
        RECT 59.310 28.950 59.480 29.120 ;
        RECT 42.770 27.370 42.940 27.540 ;
        RECT 36.810 26.550 36.980 26.720 ;
        RECT 33.760 26.140 33.930 26.310 ;
        RECT 35.400 26.140 35.570 26.310 ;
        RECT 36.310 26.140 36.480 26.310 ;
        RECT 37.920 26.180 38.090 26.350 ;
        RECT 40.610 26.890 40.780 27.060 ;
        RECT 49.030 27.810 49.200 27.980 ;
        RECT 49.950 27.810 50.120 27.980 ;
        RECT 51.580 27.720 51.750 27.890 ;
        RECT 58.870 28.090 59.040 28.260 ;
        RECT 60.920 28.990 61.090 29.160 ;
        RECT 63.610 29.700 63.780 29.870 ;
        RECT 72.030 30.620 72.200 30.790 ;
        RECT 72.950 30.620 73.120 30.790 ;
        RECT 74.580 30.530 74.750 30.700 ;
        RECT 81.870 30.820 82.040 30.990 ;
        RECT 71.520 30.180 71.690 30.350 ;
        RECT 65.560 29.360 65.730 29.530 ;
        RECT 62.510 28.950 62.680 29.120 ;
        RECT 64.150 28.950 64.320 29.120 ;
        RECT 65.060 28.950 65.230 29.120 ;
        RECT 48.520 27.370 48.690 27.540 ;
        RECT 42.560 26.550 42.730 26.720 ;
        RECT 39.510 26.140 39.680 26.310 ;
        RECT 41.150 26.140 41.320 26.310 ;
        RECT 42.060 26.140 42.230 26.310 ;
        RECT 43.670 26.180 43.840 26.350 ;
        RECT 46.360 26.890 46.530 27.060 ;
        RECT 54.780 27.810 54.950 27.980 ;
        RECT 55.700 27.810 55.870 27.980 ;
        RECT 57.330 27.720 57.500 27.890 ;
        RECT 64.620 28.090 64.790 28.260 ;
        RECT 66.670 28.990 66.840 29.160 ;
        RECT 69.360 29.700 69.530 29.870 ;
        RECT 77.780 30.620 77.950 30.790 ;
        RECT 78.700 30.620 78.870 30.790 ;
        RECT 80.330 30.530 80.500 30.700 ;
        RECT 87.620 30.820 87.790 30.990 ;
        RECT 77.270 30.180 77.440 30.350 ;
        RECT 71.310 29.360 71.480 29.530 ;
        RECT 68.260 28.950 68.430 29.120 ;
        RECT 69.900 28.950 70.070 29.120 ;
        RECT 70.810 28.950 70.980 29.120 ;
        RECT 54.270 27.370 54.440 27.540 ;
        RECT 48.310 26.550 48.480 26.720 ;
        RECT 45.260 26.140 45.430 26.310 ;
        RECT 46.900 26.140 47.070 26.310 ;
        RECT 47.810 26.140 47.980 26.310 ;
        RECT 49.420 26.180 49.590 26.350 ;
        RECT 52.110 26.890 52.280 27.060 ;
        RECT 60.530 27.810 60.700 27.980 ;
        RECT 61.450 27.810 61.620 27.980 ;
        RECT 63.080 27.720 63.250 27.890 ;
        RECT 70.370 28.090 70.540 28.260 ;
        RECT 72.420 28.990 72.590 29.160 ;
        RECT 75.110 29.700 75.280 29.870 ;
        RECT 83.530 30.620 83.700 30.790 ;
        RECT 84.450 30.620 84.620 30.790 ;
        RECT 86.080 30.530 86.250 30.700 ;
        RECT 93.370 30.820 93.540 30.990 ;
        RECT 83.020 30.180 83.190 30.350 ;
        RECT 77.060 29.360 77.230 29.530 ;
        RECT 74.010 28.950 74.180 29.120 ;
        RECT 75.650 28.950 75.820 29.120 ;
        RECT 76.560 28.950 76.730 29.120 ;
        RECT 60.020 27.370 60.190 27.540 ;
        RECT 54.060 26.550 54.230 26.720 ;
        RECT 51.010 26.140 51.180 26.310 ;
        RECT 52.650 26.140 52.820 26.310 ;
        RECT 53.560 26.140 53.730 26.310 ;
        RECT 55.170 26.180 55.340 26.350 ;
        RECT 57.860 26.890 58.030 27.060 ;
        RECT 66.280 27.810 66.450 27.980 ;
        RECT 67.200 27.810 67.370 27.980 ;
        RECT 68.830 27.720 69.000 27.890 ;
        RECT 76.120 28.090 76.290 28.260 ;
        RECT 78.170 28.990 78.340 29.160 ;
        RECT 80.860 29.700 81.030 29.870 ;
        RECT 89.280 30.620 89.450 30.790 ;
        RECT 90.200 30.620 90.370 30.790 ;
        RECT 91.830 30.530 92.000 30.700 ;
        RECT 88.770 30.180 88.940 30.350 ;
        RECT 82.810 29.360 82.980 29.530 ;
        RECT 79.760 28.950 79.930 29.120 ;
        RECT 81.400 28.950 81.570 29.120 ;
        RECT 82.310 28.950 82.480 29.120 ;
        RECT 65.770 27.370 65.940 27.540 ;
        RECT 59.810 26.550 59.980 26.720 ;
        RECT 56.760 26.140 56.930 26.310 ;
        RECT 58.400 26.140 58.570 26.310 ;
        RECT 59.310 26.140 59.480 26.310 ;
        RECT 60.920 26.180 61.090 26.350 ;
        RECT 63.610 26.890 63.780 27.060 ;
        RECT 72.030 27.810 72.200 27.980 ;
        RECT 72.950 27.810 73.120 27.980 ;
        RECT 74.580 27.720 74.750 27.890 ;
        RECT 81.870 28.090 82.040 28.260 ;
        RECT 83.920 28.990 84.090 29.160 ;
        RECT 86.610 29.700 86.780 29.870 ;
        RECT 88.560 29.360 88.730 29.530 ;
        RECT 85.510 28.950 85.680 29.120 ;
        RECT 87.150 28.950 87.320 29.120 ;
        RECT 88.060 28.950 88.230 29.120 ;
        RECT 71.520 27.370 71.690 27.540 ;
        RECT 65.560 26.550 65.730 26.720 ;
        RECT 62.510 26.140 62.680 26.310 ;
        RECT 64.150 26.140 64.320 26.310 ;
        RECT 65.060 26.140 65.230 26.310 ;
        RECT 66.670 26.180 66.840 26.350 ;
        RECT 69.360 26.890 69.530 27.060 ;
        RECT 77.780 27.810 77.950 27.980 ;
        RECT 78.700 27.810 78.870 27.980 ;
        RECT 80.330 27.720 80.500 27.890 ;
        RECT 87.620 28.090 87.790 28.260 ;
        RECT 89.670 28.990 89.840 29.160 ;
        RECT 92.360 29.700 92.530 29.870 ;
        RECT 94.310 29.360 94.480 29.530 ;
        RECT 91.260 28.950 91.430 29.120 ;
        RECT 92.900 28.950 93.070 29.120 ;
        RECT 93.810 28.950 93.980 29.120 ;
        RECT 77.270 27.370 77.440 27.540 ;
        RECT 71.310 26.550 71.480 26.720 ;
        RECT 68.260 26.140 68.430 26.310 ;
        RECT 69.900 26.140 70.070 26.310 ;
        RECT 70.810 26.140 70.980 26.310 ;
        RECT 72.420 26.180 72.590 26.350 ;
        RECT 75.110 26.890 75.280 27.060 ;
        RECT 83.530 27.810 83.700 27.980 ;
        RECT 84.450 27.810 84.620 27.980 ;
        RECT 86.080 27.720 86.250 27.890 ;
        RECT 83.020 27.370 83.190 27.540 ;
        RECT 77.060 26.550 77.230 26.720 ;
        RECT 74.010 26.140 74.180 26.310 ;
        RECT 75.650 26.140 75.820 26.310 ;
        RECT 76.560 26.140 76.730 26.310 ;
        RECT 78.170 26.180 78.340 26.350 ;
        RECT 80.860 26.890 81.030 27.060 ;
        RECT 89.280 27.810 89.450 27.980 ;
        RECT 90.200 27.810 90.370 27.980 ;
        RECT 91.830 27.720 92.000 27.890 ;
        RECT 88.770 27.370 88.940 27.540 ;
        RECT 82.810 26.550 82.980 26.720 ;
        RECT 79.760 26.140 79.930 26.310 ;
        RECT 81.400 26.140 81.570 26.310 ;
        RECT 82.310 26.140 82.480 26.310 ;
        RECT 83.920 26.180 84.090 26.350 ;
        RECT 86.610 26.890 86.780 27.060 ;
        RECT 88.560 26.550 88.730 26.720 ;
        RECT 85.510 26.140 85.680 26.310 ;
        RECT 87.150 26.140 87.320 26.310 ;
        RECT 88.060 26.140 88.230 26.310 ;
        RECT 89.670 26.180 89.840 26.350 ;
        RECT 92.360 26.890 92.530 27.060 ;
        RECT 94.310 26.550 94.480 26.720 ;
        RECT 91.260 26.140 91.430 26.310 ;
        RECT 92.900 26.140 93.070 26.310 ;
        RECT 93.810 26.140 93.980 26.310 ;
        RECT 7.120 25.600 7.290 25.770 ;
        RECT 3.030 25.400 3.200 25.570 ;
        RECT 3.950 25.400 4.120 25.570 ;
        RECT 5.580 25.310 5.750 25.480 ;
        RECT 12.870 25.600 13.040 25.770 ;
        RECT 2.520 24.960 2.690 25.130 ;
        RECT 8.780 25.400 8.950 25.570 ;
        RECT 9.700 25.400 9.870 25.570 ;
        RECT 11.330 25.310 11.500 25.480 ;
        RECT 18.620 25.600 18.790 25.770 ;
        RECT 8.270 24.960 8.440 25.130 ;
        RECT 3.420 23.770 3.590 23.940 ;
        RECT 6.110 24.480 6.280 24.650 ;
        RECT 14.530 25.400 14.700 25.570 ;
        RECT 15.450 25.400 15.620 25.570 ;
        RECT 17.080 25.310 17.250 25.480 ;
        RECT 24.370 25.600 24.540 25.770 ;
        RECT 14.020 24.960 14.190 25.130 ;
        RECT 8.060 24.140 8.230 24.310 ;
        RECT 5.010 23.730 5.180 23.900 ;
        RECT 6.650 23.730 6.820 23.900 ;
        RECT 7.560 23.730 7.730 23.900 ;
        RECT 9.170 23.770 9.340 23.940 ;
        RECT 11.860 24.480 12.030 24.650 ;
        RECT 20.280 25.400 20.450 25.570 ;
        RECT 21.200 25.400 21.370 25.570 ;
        RECT 22.830 25.310 23.000 25.480 ;
        RECT 30.120 25.600 30.290 25.770 ;
        RECT 19.770 24.960 19.940 25.130 ;
        RECT 13.810 24.140 13.980 24.310 ;
        RECT 10.760 23.730 10.930 23.900 ;
        RECT 12.400 23.730 12.570 23.900 ;
        RECT 13.310 23.730 13.480 23.900 ;
        RECT 14.920 23.770 15.090 23.940 ;
        RECT 17.610 24.480 17.780 24.650 ;
        RECT 26.030 25.400 26.200 25.570 ;
        RECT 26.950 25.400 27.120 25.570 ;
        RECT 28.580 25.310 28.750 25.480 ;
        RECT 35.870 25.600 36.040 25.770 ;
        RECT 25.520 24.960 25.690 25.130 ;
        RECT 19.560 24.140 19.730 24.310 ;
        RECT 16.510 23.730 16.680 23.900 ;
        RECT 18.150 23.730 18.320 23.900 ;
        RECT 19.060 23.730 19.230 23.900 ;
        RECT 20.670 23.770 20.840 23.940 ;
        RECT 23.360 24.480 23.530 24.650 ;
        RECT 31.780 25.400 31.950 25.570 ;
        RECT 32.700 25.400 32.870 25.570 ;
        RECT 34.330 25.310 34.500 25.480 ;
        RECT 41.620 25.600 41.790 25.770 ;
        RECT 31.270 24.960 31.440 25.130 ;
        RECT 25.310 24.140 25.480 24.310 ;
        RECT 22.260 23.730 22.430 23.900 ;
        RECT 23.900 23.730 24.070 23.900 ;
        RECT 24.810 23.730 24.980 23.900 ;
        RECT 26.420 23.770 26.590 23.940 ;
        RECT 29.110 24.480 29.280 24.650 ;
        RECT 37.530 25.400 37.700 25.570 ;
        RECT 38.450 25.400 38.620 25.570 ;
        RECT 40.080 25.310 40.250 25.480 ;
        RECT 47.370 25.600 47.540 25.770 ;
        RECT 37.020 24.960 37.190 25.130 ;
        RECT 31.060 24.140 31.230 24.310 ;
        RECT 28.010 23.730 28.180 23.900 ;
        RECT 29.650 23.730 29.820 23.900 ;
        RECT 30.560 23.730 30.730 23.900 ;
        RECT 32.170 23.770 32.340 23.940 ;
        RECT 34.860 24.480 35.030 24.650 ;
        RECT 43.280 25.400 43.450 25.570 ;
        RECT 44.200 25.400 44.370 25.570 ;
        RECT 45.830 25.310 46.000 25.480 ;
        RECT 53.120 25.600 53.290 25.770 ;
        RECT 42.770 24.960 42.940 25.130 ;
        RECT 36.810 24.140 36.980 24.310 ;
        RECT 33.760 23.730 33.930 23.900 ;
        RECT 35.400 23.730 35.570 23.900 ;
        RECT 36.310 23.730 36.480 23.900 ;
        RECT 37.920 23.770 38.090 23.940 ;
        RECT 40.610 24.480 40.780 24.650 ;
        RECT 49.030 25.400 49.200 25.570 ;
        RECT 49.950 25.400 50.120 25.570 ;
        RECT 51.580 25.310 51.750 25.480 ;
        RECT 58.870 25.600 59.040 25.770 ;
        RECT 48.520 24.960 48.690 25.130 ;
        RECT 42.560 24.140 42.730 24.310 ;
        RECT 39.510 23.730 39.680 23.900 ;
        RECT 41.150 23.730 41.320 23.900 ;
        RECT 42.060 23.730 42.230 23.900 ;
        RECT 43.670 23.770 43.840 23.940 ;
        RECT 46.360 24.480 46.530 24.650 ;
        RECT 54.780 25.400 54.950 25.570 ;
        RECT 55.700 25.400 55.870 25.570 ;
        RECT 57.330 25.310 57.500 25.480 ;
        RECT 64.620 25.600 64.790 25.770 ;
        RECT 54.270 24.960 54.440 25.130 ;
        RECT 48.310 24.140 48.480 24.310 ;
        RECT 45.260 23.730 45.430 23.900 ;
        RECT 46.900 23.730 47.070 23.900 ;
        RECT 47.810 23.730 47.980 23.900 ;
        RECT 49.420 23.770 49.590 23.940 ;
        RECT 52.110 24.480 52.280 24.650 ;
        RECT 60.530 25.400 60.700 25.570 ;
        RECT 61.450 25.400 61.620 25.570 ;
        RECT 63.080 25.310 63.250 25.480 ;
        RECT 70.370 25.600 70.540 25.770 ;
        RECT 60.020 24.960 60.190 25.130 ;
        RECT 54.060 24.140 54.230 24.310 ;
        RECT 51.010 23.730 51.180 23.900 ;
        RECT 52.650 23.730 52.820 23.900 ;
        RECT 53.560 23.730 53.730 23.900 ;
        RECT 55.170 23.770 55.340 23.940 ;
        RECT 57.860 24.480 58.030 24.650 ;
        RECT 66.280 25.400 66.450 25.570 ;
        RECT 67.200 25.400 67.370 25.570 ;
        RECT 68.830 25.310 69.000 25.480 ;
        RECT 76.120 25.600 76.290 25.770 ;
        RECT 65.770 24.960 65.940 25.130 ;
        RECT 59.810 24.140 59.980 24.310 ;
        RECT 56.760 23.730 56.930 23.900 ;
        RECT 58.400 23.730 58.570 23.900 ;
        RECT 59.310 23.730 59.480 23.900 ;
        RECT 60.920 23.770 61.090 23.940 ;
        RECT 63.610 24.480 63.780 24.650 ;
        RECT 72.030 25.400 72.200 25.570 ;
        RECT 72.950 25.400 73.120 25.570 ;
        RECT 74.580 25.310 74.750 25.480 ;
        RECT 81.870 25.600 82.040 25.770 ;
        RECT 71.520 24.960 71.690 25.130 ;
        RECT 65.560 24.140 65.730 24.310 ;
        RECT 62.510 23.730 62.680 23.900 ;
        RECT 64.150 23.730 64.320 23.900 ;
        RECT 65.060 23.730 65.230 23.900 ;
        RECT 66.670 23.770 66.840 23.940 ;
        RECT 69.360 24.480 69.530 24.650 ;
        RECT 77.780 25.400 77.950 25.570 ;
        RECT 78.700 25.400 78.870 25.570 ;
        RECT 80.330 25.310 80.500 25.480 ;
        RECT 87.620 25.600 87.790 25.770 ;
        RECT 77.270 24.960 77.440 25.130 ;
        RECT 71.310 24.140 71.480 24.310 ;
        RECT 68.260 23.730 68.430 23.900 ;
        RECT 69.900 23.730 70.070 23.900 ;
        RECT 70.810 23.730 70.980 23.900 ;
        RECT 72.420 23.770 72.590 23.940 ;
        RECT 75.110 24.480 75.280 24.650 ;
        RECT 83.530 25.400 83.700 25.570 ;
        RECT 84.450 25.400 84.620 25.570 ;
        RECT 86.080 25.310 86.250 25.480 ;
        RECT 93.370 25.600 93.540 25.770 ;
        RECT 83.020 24.960 83.190 25.130 ;
        RECT 77.060 24.140 77.230 24.310 ;
        RECT 74.010 23.730 74.180 23.900 ;
        RECT 75.650 23.730 75.820 23.900 ;
        RECT 76.560 23.730 76.730 23.900 ;
        RECT 78.170 23.770 78.340 23.940 ;
        RECT 80.860 24.480 81.030 24.650 ;
        RECT 89.280 25.400 89.450 25.570 ;
        RECT 90.200 25.400 90.370 25.570 ;
        RECT 91.830 25.310 92.000 25.480 ;
        RECT 88.770 24.960 88.940 25.130 ;
        RECT 82.810 24.140 82.980 24.310 ;
        RECT 79.760 23.730 79.930 23.900 ;
        RECT 81.400 23.730 81.570 23.900 ;
        RECT 82.310 23.730 82.480 23.900 ;
        RECT 83.920 23.770 84.090 23.940 ;
        RECT 86.610 24.480 86.780 24.650 ;
        RECT 88.560 24.140 88.730 24.310 ;
        RECT 85.510 23.730 85.680 23.900 ;
        RECT 87.150 23.730 87.320 23.900 ;
        RECT 88.060 23.730 88.230 23.900 ;
        RECT 89.670 23.770 89.840 23.940 ;
        RECT 92.360 24.480 92.530 24.650 ;
        RECT 94.310 24.140 94.480 24.310 ;
        RECT 91.260 23.730 91.430 23.900 ;
        RECT 92.900 23.730 93.070 23.900 ;
        RECT 93.810 23.730 93.980 23.900 ;
        RECT 7.120 23.190 7.290 23.360 ;
        RECT 3.030 22.990 3.200 23.160 ;
        RECT 3.950 22.990 4.120 23.160 ;
        RECT 5.580 22.900 5.750 23.070 ;
        RECT 12.870 23.190 13.040 23.360 ;
        RECT 2.520 22.550 2.690 22.720 ;
        RECT 8.780 22.990 8.950 23.160 ;
        RECT 9.700 22.990 9.870 23.160 ;
        RECT 11.330 22.900 11.500 23.070 ;
        RECT 18.620 23.190 18.790 23.360 ;
        RECT 8.270 22.550 8.440 22.720 ;
        RECT 3.420 21.360 3.590 21.530 ;
        RECT 6.110 22.070 6.280 22.240 ;
        RECT 14.530 22.990 14.700 23.160 ;
        RECT 15.450 22.990 15.620 23.160 ;
        RECT 17.080 22.900 17.250 23.070 ;
        RECT 24.370 23.190 24.540 23.360 ;
        RECT 14.020 22.550 14.190 22.720 ;
        RECT 8.060 21.730 8.230 21.900 ;
        RECT 5.010 21.320 5.180 21.490 ;
        RECT 6.650 21.320 6.820 21.490 ;
        RECT 7.560 21.320 7.730 21.490 ;
        RECT 9.170 21.360 9.340 21.530 ;
        RECT 11.860 22.070 12.030 22.240 ;
        RECT 20.280 22.990 20.450 23.160 ;
        RECT 21.200 22.990 21.370 23.160 ;
        RECT 22.830 22.900 23.000 23.070 ;
        RECT 30.120 23.190 30.290 23.360 ;
        RECT 19.770 22.550 19.940 22.720 ;
        RECT 13.810 21.730 13.980 21.900 ;
        RECT 10.760 21.320 10.930 21.490 ;
        RECT 12.400 21.320 12.570 21.490 ;
        RECT 13.310 21.320 13.480 21.490 ;
        RECT 14.920 21.360 15.090 21.530 ;
        RECT 17.610 22.070 17.780 22.240 ;
        RECT 26.030 22.990 26.200 23.160 ;
        RECT 26.950 22.990 27.120 23.160 ;
        RECT 28.580 22.900 28.750 23.070 ;
        RECT 35.870 23.190 36.040 23.360 ;
        RECT 25.520 22.550 25.690 22.720 ;
        RECT 19.560 21.730 19.730 21.900 ;
        RECT 16.510 21.320 16.680 21.490 ;
        RECT 18.150 21.320 18.320 21.490 ;
        RECT 19.060 21.320 19.230 21.490 ;
        RECT 20.670 21.360 20.840 21.530 ;
        RECT 23.360 22.070 23.530 22.240 ;
        RECT 31.780 22.990 31.950 23.160 ;
        RECT 32.700 22.990 32.870 23.160 ;
        RECT 34.330 22.900 34.500 23.070 ;
        RECT 41.620 23.190 41.790 23.360 ;
        RECT 31.270 22.550 31.440 22.720 ;
        RECT 25.310 21.730 25.480 21.900 ;
        RECT 22.260 21.320 22.430 21.490 ;
        RECT 23.900 21.320 24.070 21.490 ;
        RECT 24.810 21.320 24.980 21.490 ;
        RECT 26.420 21.360 26.590 21.530 ;
        RECT 29.110 22.070 29.280 22.240 ;
        RECT 37.530 22.990 37.700 23.160 ;
        RECT 38.450 22.990 38.620 23.160 ;
        RECT 40.080 22.900 40.250 23.070 ;
        RECT 47.370 23.190 47.540 23.360 ;
        RECT 37.020 22.550 37.190 22.720 ;
        RECT 31.060 21.730 31.230 21.900 ;
        RECT 28.010 21.320 28.180 21.490 ;
        RECT 29.650 21.320 29.820 21.490 ;
        RECT 30.560 21.320 30.730 21.490 ;
        RECT 32.170 21.360 32.340 21.530 ;
        RECT 34.860 22.070 35.030 22.240 ;
        RECT 43.280 22.990 43.450 23.160 ;
        RECT 44.200 22.990 44.370 23.160 ;
        RECT 45.830 22.900 46.000 23.070 ;
        RECT 53.120 23.190 53.290 23.360 ;
        RECT 42.770 22.550 42.940 22.720 ;
        RECT 36.810 21.730 36.980 21.900 ;
        RECT 33.760 21.320 33.930 21.490 ;
        RECT 35.400 21.320 35.570 21.490 ;
        RECT 36.310 21.320 36.480 21.490 ;
        RECT 37.920 21.360 38.090 21.530 ;
        RECT 40.610 22.070 40.780 22.240 ;
        RECT 49.030 22.990 49.200 23.160 ;
        RECT 49.950 22.990 50.120 23.160 ;
        RECT 51.580 22.900 51.750 23.070 ;
        RECT 58.870 23.190 59.040 23.360 ;
        RECT 48.520 22.550 48.690 22.720 ;
        RECT 42.560 21.730 42.730 21.900 ;
        RECT 39.510 21.320 39.680 21.490 ;
        RECT 41.150 21.320 41.320 21.490 ;
        RECT 42.060 21.320 42.230 21.490 ;
        RECT 43.670 21.360 43.840 21.530 ;
        RECT 46.360 22.070 46.530 22.240 ;
        RECT 54.780 22.990 54.950 23.160 ;
        RECT 55.700 22.990 55.870 23.160 ;
        RECT 57.330 22.900 57.500 23.070 ;
        RECT 64.620 23.190 64.790 23.360 ;
        RECT 54.270 22.550 54.440 22.720 ;
        RECT 48.310 21.730 48.480 21.900 ;
        RECT 45.260 21.320 45.430 21.490 ;
        RECT 46.900 21.320 47.070 21.490 ;
        RECT 47.810 21.320 47.980 21.490 ;
        RECT 49.420 21.360 49.590 21.530 ;
        RECT 52.110 22.070 52.280 22.240 ;
        RECT 60.530 22.990 60.700 23.160 ;
        RECT 61.450 22.990 61.620 23.160 ;
        RECT 63.080 22.900 63.250 23.070 ;
        RECT 70.370 23.190 70.540 23.360 ;
        RECT 60.020 22.550 60.190 22.720 ;
        RECT 54.060 21.730 54.230 21.900 ;
        RECT 51.010 21.320 51.180 21.490 ;
        RECT 52.650 21.320 52.820 21.490 ;
        RECT 53.560 21.320 53.730 21.490 ;
        RECT 55.170 21.360 55.340 21.530 ;
        RECT 57.860 22.070 58.030 22.240 ;
        RECT 66.280 22.990 66.450 23.160 ;
        RECT 67.200 22.990 67.370 23.160 ;
        RECT 68.830 22.900 69.000 23.070 ;
        RECT 76.120 23.190 76.290 23.360 ;
        RECT 65.770 22.550 65.940 22.720 ;
        RECT 59.810 21.730 59.980 21.900 ;
        RECT 56.760 21.320 56.930 21.490 ;
        RECT 58.400 21.320 58.570 21.490 ;
        RECT 59.310 21.320 59.480 21.490 ;
        RECT 60.920 21.360 61.090 21.530 ;
        RECT 63.610 22.070 63.780 22.240 ;
        RECT 72.030 22.990 72.200 23.160 ;
        RECT 72.950 22.990 73.120 23.160 ;
        RECT 74.580 22.900 74.750 23.070 ;
        RECT 81.870 23.190 82.040 23.360 ;
        RECT 71.520 22.550 71.690 22.720 ;
        RECT 65.560 21.730 65.730 21.900 ;
        RECT 62.510 21.320 62.680 21.490 ;
        RECT 64.150 21.320 64.320 21.490 ;
        RECT 65.060 21.320 65.230 21.490 ;
        RECT 66.670 21.360 66.840 21.530 ;
        RECT 69.360 22.070 69.530 22.240 ;
        RECT 77.780 22.990 77.950 23.160 ;
        RECT 78.700 22.990 78.870 23.160 ;
        RECT 80.330 22.900 80.500 23.070 ;
        RECT 87.620 23.190 87.790 23.360 ;
        RECT 77.270 22.550 77.440 22.720 ;
        RECT 71.310 21.730 71.480 21.900 ;
        RECT 68.260 21.320 68.430 21.490 ;
        RECT 69.900 21.320 70.070 21.490 ;
        RECT 70.810 21.320 70.980 21.490 ;
        RECT 72.420 21.360 72.590 21.530 ;
        RECT 75.110 22.070 75.280 22.240 ;
        RECT 83.530 22.990 83.700 23.160 ;
        RECT 84.450 22.990 84.620 23.160 ;
        RECT 86.080 22.900 86.250 23.070 ;
        RECT 93.370 23.190 93.540 23.360 ;
        RECT 83.020 22.550 83.190 22.720 ;
        RECT 77.060 21.730 77.230 21.900 ;
        RECT 74.010 21.320 74.180 21.490 ;
        RECT 75.650 21.320 75.820 21.490 ;
        RECT 76.560 21.320 76.730 21.490 ;
        RECT 78.170 21.360 78.340 21.530 ;
        RECT 80.860 22.070 81.030 22.240 ;
        RECT 89.280 22.990 89.450 23.160 ;
        RECT 90.200 22.990 90.370 23.160 ;
        RECT 91.830 22.900 92.000 23.070 ;
        RECT 88.770 22.550 88.940 22.720 ;
        RECT 82.810 21.730 82.980 21.900 ;
        RECT 79.760 21.320 79.930 21.490 ;
        RECT 81.400 21.320 81.570 21.490 ;
        RECT 82.310 21.320 82.480 21.490 ;
        RECT 83.920 21.360 84.090 21.530 ;
        RECT 86.610 22.070 86.780 22.240 ;
        RECT 88.560 21.730 88.730 21.900 ;
        RECT 85.510 21.320 85.680 21.490 ;
        RECT 87.150 21.320 87.320 21.490 ;
        RECT 88.060 21.320 88.230 21.490 ;
        RECT 89.670 21.360 89.840 21.530 ;
        RECT 92.360 22.070 92.530 22.240 ;
        RECT 94.310 21.730 94.480 21.900 ;
        RECT 91.260 21.320 91.430 21.490 ;
        RECT 92.900 21.320 93.070 21.490 ;
        RECT 93.810 21.320 93.980 21.490 ;
        RECT 7.120 20.780 7.290 20.950 ;
        RECT 3.030 20.580 3.200 20.750 ;
        RECT 3.950 20.580 4.120 20.750 ;
        RECT 5.580 20.490 5.750 20.660 ;
        RECT 12.870 20.780 13.040 20.950 ;
        RECT 2.520 20.140 2.690 20.310 ;
        RECT 8.780 20.580 8.950 20.750 ;
        RECT 9.700 20.580 9.870 20.750 ;
        RECT 11.330 20.490 11.500 20.660 ;
        RECT 18.620 20.780 18.790 20.950 ;
        RECT 8.270 20.140 8.440 20.310 ;
        RECT 3.420 18.950 3.590 19.120 ;
        RECT 6.110 19.660 6.280 19.830 ;
        RECT 14.530 20.580 14.700 20.750 ;
        RECT 15.450 20.580 15.620 20.750 ;
        RECT 17.080 20.490 17.250 20.660 ;
        RECT 24.370 20.780 24.540 20.950 ;
        RECT 14.020 20.140 14.190 20.310 ;
        RECT 8.060 19.320 8.230 19.490 ;
        RECT 5.010 18.910 5.180 19.080 ;
        RECT 6.650 18.910 6.820 19.080 ;
        RECT 7.560 18.910 7.730 19.080 ;
        RECT 9.170 18.950 9.340 19.120 ;
        RECT 11.860 19.660 12.030 19.830 ;
        RECT 20.280 20.580 20.450 20.750 ;
        RECT 21.200 20.580 21.370 20.750 ;
        RECT 22.830 20.490 23.000 20.660 ;
        RECT 30.120 20.780 30.290 20.950 ;
        RECT 19.770 20.140 19.940 20.310 ;
        RECT 13.810 19.320 13.980 19.490 ;
        RECT 10.760 18.910 10.930 19.080 ;
        RECT 12.400 18.910 12.570 19.080 ;
        RECT 13.310 18.910 13.480 19.080 ;
        RECT 14.920 18.950 15.090 19.120 ;
        RECT 17.610 19.660 17.780 19.830 ;
        RECT 26.030 20.580 26.200 20.750 ;
        RECT 26.950 20.580 27.120 20.750 ;
        RECT 28.580 20.490 28.750 20.660 ;
        RECT 35.870 20.780 36.040 20.950 ;
        RECT 25.520 20.140 25.690 20.310 ;
        RECT 19.560 19.320 19.730 19.490 ;
        RECT 16.510 18.910 16.680 19.080 ;
        RECT 18.150 18.910 18.320 19.080 ;
        RECT 19.060 18.910 19.230 19.080 ;
        RECT 20.670 18.950 20.840 19.120 ;
        RECT 23.360 19.660 23.530 19.830 ;
        RECT 31.780 20.580 31.950 20.750 ;
        RECT 32.700 20.580 32.870 20.750 ;
        RECT 34.330 20.490 34.500 20.660 ;
        RECT 41.620 20.780 41.790 20.950 ;
        RECT 31.270 20.140 31.440 20.310 ;
        RECT 25.310 19.320 25.480 19.490 ;
        RECT 22.260 18.910 22.430 19.080 ;
        RECT 23.900 18.910 24.070 19.080 ;
        RECT 24.810 18.910 24.980 19.080 ;
        RECT 26.420 18.950 26.590 19.120 ;
        RECT 29.110 19.660 29.280 19.830 ;
        RECT 37.530 20.580 37.700 20.750 ;
        RECT 38.450 20.580 38.620 20.750 ;
        RECT 40.080 20.490 40.250 20.660 ;
        RECT 47.370 20.780 47.540 20.950 ;
        RECT 37.020 20.140 37.190 20.310 ;
        RECT 31.060 19.320 31.230 19.490 ;
        RECT 28.010 18.910 28.180 19.080 ;
        RECT 29.650 18.910 29.820 19.080 ;
        RECT 30.560 18.910 30.730 19.080 ;
        RECT 32.170 18.950 32.340 19.120 ;
        RECT 34.860 19.660 35.030 19.830 ;
        RECT 43.280 20.580 43.450 20.750 ;
        RECT 44.200 20.580 44.370 20.750 ;
        RECT 45.830 20.490 46.000 20.660 ;
        RECT 53.120 20.780 53.290 20.950 ;
        RECT 42.770 20.140 42.940 20.310 ;
        RECT 36.810 19.320 36.980 19.490 ;
        RECT 33.760 18.910 33.930 19.080 ;
        RECT 35.400 18.910 35.570 19.080 ;
        RECT 36.310 18.910 36.480 19.080 ;
        RECT 37.920 18.950 38.090 19.120 ;
        RECT 40.610 19.660 40.780 19.830 ;
        RECT 49.030 20.580 49.200 20.750 ;
        RECT 49.950 20.580 50.120 20.750 ;
        RECT 51.580 20.490 51.750 20.660 ;
        RECT 58.870 20.780 59.040 20.950 ;
        RECT 48.520 20.140 48.690 20.310 ;
        RECT 42.560 19.320 42.730 19.490 ;
        RECT 39.510 18.910 39.680 19.080 ;
        RECT 41.150 18.910 41.320 19.080 ;
        RECT 42.060 18.910 42.230 19.080 ;
        RECT 43.670 18.950 43.840 19.120 ;
        RECT 46.360 19.660 46.530 19.830 ;
        RECT 54.780 20.580 54.950 20.750 ;
        RECT 55.700 20.580 55.870 20.750 ;
        RECT 57.330 20.490 57.500 20.660 ;
        RECT 64.620 20.780 64.790 20.950 ;
        RECT 54.270 20.140 54.440 20.310 ;
        RECT 48.310 19.320 48.480 19.490 ;
        RECT 45.260 18.910 45.430 19.080 ;
        RECT 46.900 18.910 47.070 19.080 ;
        RECT 47.810 18.910 47.980 19.080 ;
        RECT 49.420 18.950 49.590 19.120 ;
        RECT 52.110 19.660 52.280 19.830 ;
        RECT 60.530 20.580 60.700 20.750 ;
        RECT 61.450 20.580 61.620 20.750 ;
        RECT 63.080 20.490 63.250 20.660 ;
        RECT 70.370 20.780 70.540 20.950 ;
        RECT 60.020 20.140 60.190 20.310 ;
        RECT 54.060 19.320 54.230 19.490 ;
        RECT 51.010 18.910 51.180 19.080 ;
        RECT 52.650 18.910 52.820 19.080 ;
        RECT 53.560 18.910 53.730 19.080 ;
        RECT 55.170 18.950 55.340 19.120 ;
        RECT 57.860 19.660 58.030 19.830 ;
        RECT 66.280 20.580 66.450 20.750 ;
        RECT 67.200 20.580 67.370 20.750 ;
        RECT 68.830 20.490 69.000 20.660 ;
        RECT 76.120 20.780 76.290 20.950 ;
        RECT 65.770 20.140 65.940 20.310 ;
        RECT 59.810 19.320 59.980 19.490 ;
        RECT 56.760 18.910 56.930 19.080 ;
        RECT 58.400 18.910 58.570 19.080 ;
        RECT 59.310 18.910 59.480 19.080 ;
        RECT 60.920 18.950 61.090 19.120 ;
        RECT 63.610 19.660 63.780 19.830 ;
        RECT 72.030 20.580 72.200 20.750 ;
        RECT 72.950 20.580 73.120 20.750 ;
        RECT 74.580 20.490 74.750 20.660 ;
        RECT 81.870 20.780 82.040 20.950 ;
        RECT 71.520 20.140 71.690 20.310 ;
        RECT 65.560 19.320 65.730 19.490 ;
        RECT 62.510 18.910 62.680 19.080 ;
        RECT 64.150 18.910 64.320 19.080 ;
        RECT 65.060 18.910 65.230 19.080 ;
        RECT 66.670 18.950 66.840 19.120 ;
        RECT 69.360 19.660 69.530 19.830 ;
        RECT 77.780 20.580 77.950 20.750 ;
        RECT 78.700 20.580 78.870 20.750 ;
        RECT 80.330 20.490 80.500 20.660 ;
        RECT 87.620 20.780 87.790 20.950 ;
        RECT 77.270 20.140 77.440 20.310 ;
        RECT 71.310 19.320 71.480 19.490 ;
        RECT 68.260 18.910 68.430 19.080 ;
        RECT 69.900 18.910 70.070 19.080 ;
        RECT 70.810 18.910 70.980 19.080 ;
        RECT 72.420 18.950 72.590 19.120 ;
        RECT 75.110 19.660 75.280 19.830 ;
        RECT 83.530 20.580 83.700 20.750 ;
        RECT 84.450 20.580 84.620 20.750 ;
        RECT 86.080 20.490 86.250 20.660 ;
        RECT 93.370 20.780 93.540 20.950 ;
        RECT 83.020 20.140 83.190 20.310 ;
        RECT 77.060 19.320 77.230 19.490 ;
        RECT 74.010 18.910 74.180 19.080 ;
        RECT 75.650 18.910 75.820 19.080 ;
        RECT 76.560 18.910 76.730 19.080 ;
        RECT 78.170 18.950 78.340 19.120 ;
        RECT 80.860 19.660 81.030 19.830 ;
        RECT 89.280 20.580 89.450 20.750 ;
        RECT 90.200 20.580 90.370 20.750 ;
        RECT 91.830 20.490 92.000 20.660 ;
        RECT 88.770 20.140 88.940 20.310 ;
        RECT 82.810 19.320 82.980 19.490 ;
        RECT 79.760 18.910 79.930 19.080 ;
        RECT 81.400 18.910 81.570 19.080 ;
        RECT 82.310 18.910 82.480 19.080 ;
        RECT 83.920 18.950 84.090 19.120 ;
        RECT 86.610 19.660 86.780 19.830 ;
        RECT 88.560 19.320 88.730 19.490 ;
        RECT 85.510 18.910 85.680 19.080 ;
        RECT 87.150 18.910 87.320 19.080 ;
        RECT 88.060 18.910 88.230 19.080 ;
        RECT 89.670 18.950 89.840 19.120 ;
        RECT 92.360 19.660 92.530 19.830 ;
        RECT 94.310 19.320 94.480 19.490 ;
        RECT 91.260 18.910 91.430 19.080 ;
        RECT 92.900 18.910 93.070 19.080 ;
        RECT 93.810 18.910 93.980 19.080 ;
        RECT 7.120 18.370 7.290 18.540 ;
        RECT 3.030 18.170 3.200 18.340 ;
        RECT 3.950 18.170 4.120 18.340 ;
        RECT 5.580 18.080 5.750 18.250 ;
        RECT 12.870 18.370 13.040 18.540 ;
        RECT 2.520 17.730 2.690 17.900 ;
        RECT 8.780 18.170 8.950 18.340 ;
        RECT 9.700 18.170 9.870 18.340 ;
        RECT 11.330 18.080 11.500 18.250 ;
        RECT 18.620 18.370 18.790 18.540 ;
        RECT 8.270 17.730 8.440 17.900 ;
        RECT 3.420 16.540 3.590 16.710 ;
        RECT 6.110 17.250 6.280 17.420 ;
        RECT 14.530 18.170 14.700 18.340 ;
        RECT 15.450 18.170 15.620 18.340 ;
        RECT 17.080 18.080 17.250 18.250 ;
        RECT 24.370 18.370 24.540 18.540 ;
        RECT 14.020 17.730 14.190 17.900 ;
        RECT 8.060 16.910 8.230 17.080 ;
        RECT 5.010 16.500 5.180 16.670 ;
        RECT 6.650 16.500 6.820 16.670 ;
        RECT 7.560 16.500 7.730 16.670 ;
        RECT 9.170 16.540 9.340 16.710 ;
        RECT 11.860 17.250 12.030 17.420 ;
        RECT 20.280 18.170 20.450 18.340 ;
        RECT 21.200 18.170 21.370 18.340 ;
        RECT 22.830 18.080 23.000 18.250 ;
        RECT 30.120 18.370 30.290 18.540 ;
        RECT 19.770 17.730 19.940 17.900 ;
        RECT 13.810 16.910 13.980 17.080 ;
        RECT 10.760 16.500 10.930 16.670 ;
        RECT 12.400 16.500 12.570 16.670 ;
        RECT 13.310 16.500 13.480 16.670 ;
        RECT 14.920 16.540 15.090 16.710 ;
        RECT 17.610 17.250 17.780 17.420 ;
        RECT 26.030 18.170 26.200 18.340 ;
        RECT 26.950 18.170 27.120 18.340 ;
        RECT 28.580 18.080 28.750 18.250 ;
        RECT 35.870 18.370 36.040 18.540 ;
        RECT 25.520 17.730 25.690 17.900 ;
        RECT 19.560 16.910 19.730 17.080 ;
        RECT 16.510 16.500 16.680 16.670 ;
        RECT 18.150 16.500 18.320 16.670 ;
        RECT 19.060 16.500 19.230 16.670 ;
        RECT 20.670 16.540 20.840 16.710 ;
        RECT 23.360 17.250 23.530 17.420 ;
        RECT 31.780 18.170 31.950 18.340 ;
        RECT 32.700 18.170 32.870 18.340 ;
        RECT 34.330 18.080 34.500 18.250 ;
        RECT 41.620 18.370 41.790 18.540 ;
        RECT 31.270 17.730 31.440 17.900 ;
        RECT 25.310 16.910 25.480 17.080 ;
        RECT 22.260 16.500 22.430 16.670 ;
        RECT 23.900 16.500 24.070 16.670 ;
        RECT 24.810 16.500 24.980 16.670 ;
        RECT 26.420 16.540 26.590 16.710 ;
        RECT 29.110 17.250 29.280 17.420 ;
        RECT 37.530 18.170 37.700 18.340 ;
        RECT 38.450 18.170 38.620 18.340 ;
        RECT 40.080 18.080 40.250 18.250 ;
        RECT 47.370 18.370 47.540 18.540 ;
        RECT 37.020 17.730 37.190 17.900 ;
        RECT 31.060 16.910 31.230 17.080 ;
        RECT 28.010 16.500 28.180 16.670 ;
        RECT 29.650 16.500 29.820 16.670 ;
        RECT 30.560 16.500 30.730 16.670 ;
        RECT 32.170 16.540 32.340 16.710 ;
        RECT 34.860 17.250 35.030 17.420 ;
        RECT 43.280 18.170 43.450 18.340 ;
        RECT 44.200 18.170 44.370 18.340 ;
        RECT 45.830 18.080 46.000 18.250 ;
        RECT 53.120 18.370 53.290 18.540 ;
        RECT 42.770 17.730 42.940 17.900 ;
        RECT 36.810 16.910 36.980 17.080 ;
        RECT 33.760 16.500 33.930 16.670 ;
        RECT 35.400 16.500 35.570 16.670 ;
        RECT 36.310 16.500 36.480 16.670 ;
        RECT 37.920 16.540 38.090 16.710 ;
        RECT 40.610 17.250 40.780 17.420 ;
        RECT 49.030 18.170 49.200 18.340 ;
        RECT 49.950 18.170 50.120 18.340 ;
        RECT 51.580 18.080 51.750 18.250 ;
        RECT 58.870 18.370 59.040 18.540 ;
        RECT 48.520 17.730 48.690 17.900 ;
        RECT 42.560 16.910 42.730 17.080 ;
        RECT 39.510 16.500 39.680 16.670 ;
        RECT 41.150 16.500 41.320 16.670 ;
        RECT 42.060 16.500 42.230 16.670 ;
        RECT 43.670 16.540 43.840 16.710 ;
        RECT 46.360 17.250 46.530 17.420 ;
        RECT 54.780 18.170 54.950 18.340 ;
        RECT 55.700 18.170 55.870 18.340 ;
        RECT 57.330 18.080 57.500 18.250 ;
        RECT 64.620 18.370 64.790 18.540 ;
        RECT 54.270 17.730 54.440 17.900 ;
        RECT 48.310 16.910 48.480 17.080 ;
        RECT 45.260 16.500 45.430 16.670 ;
        RECT 46.900 16.500 47.070 16.670 ;
        RECT 47.810 16.500 47.980 16.670 ;
        RECT 49.420 16.540 49.590 16.710 ;
        RECT 52.110 17.250 52.280 17.420 ;
        RECT 60.530 18.170 60.700 18.340 ;
        RECT 61.450 18.170 61.620 18.340 ;
        RECT 63.080 18.080 63.250 18.250 ;
        RECT 70.370 18.370 70.540 18.540 ;
        RECT 60.020 17.730 60.190 17.900 ;
        RECT 54.060 16.910 54.230 17.080 ;
        RECT 51.010 16.500 51.180 16.670 ;
        RECT 52.650 16.500 52.820 16.670 ;
        RECT 53.560 16.500 53.730 16.670 ;
        RECT 55.170 16.540 55.340 16.710 ;
        RECT 57.860 17.250 58.030 17.420 ;
        RECT 66.280 18.170 66.450 18.340 ;
        RECT 67.200 18.170 67.370 18.340 ;
        RECT 68.830 18.080 69.000 18.250 ;
        RECT 76.120 18.370 76.290 18.540 ;
        RECT 65.770 17.730 65.940 17.900 ;
        RECT 59.810 16.910 59.980 17.080 ;
        RECT 56.760 16.500 56.930 16.670 ;
        RECT 58.400 16.500 58.570 16.670 ;
        RECT 59.310 16.500 59.480 16.670 ;
        RECT 60.920 16.540 61.090 16.710 ;
        RECT 63.610 17.250 63.780 17.420 ;
        RECT 72.030 18.170 72.200 18.340 ;
        RECT 72.950 18.170 73.120 18.340 ;
        RECT 74.580 18.080 74.750 18.250 ;
        RECT 81.870 18.370 82.040 18.540 ;
        RECT 71.520 17.730 71.690 17.900 ;
        RECT 65.560 16.910 65.730 17.080 ;
        RECT 62.510 16.500 62.680 16.670 ;
        RECT 64.150 16.500 64.320 16.670 ;
        RECT 65.060 16.500 65.230 16.670 ;
        RECT 66.670 16.540 66.840 16.710 ;
        RECT 69.360 17.250 69.530 17.420 ;
        RECT 77.780 18.170 77.950 18.340 ;
        RECT 78.700 18.170 78.870 18.340 ;
        RECT 80.330 18.080 80.500 18.250 ;
        RECT 87.620 18.370 87.790 18.540 ;
        RECT 77.270 17.730 77.440 17.900 ;
        RECT 71.310 16.910 71.480 17.080 ;
        RECT 68.260 16.500 68.430 16.670 ;
        RECT 69.900 16.500 70.070 16.670 ;
        RECT 70.810 16.500 70.980 16.670 ;
        RECT 72.420 16.540 72.590 16.710 ;
        RECT 75.110 17.250 75.280 17.420 ;
        RECT 83.530 18.170 83.700 18.340 ;
        RECT 84.450 18.170 84.620 18.340 ;
        RECT 86.080 18.080 86.250 18.250 ;
        RECT 93.370 18.370 93.540 18.540 ;
        RECT 83.020 17.730 83.190 17.900 ;
        RECT 77.060 16.910 77.230 17.080 ;
        RECT 74.010 16.500 74.180 16.670 ;
        RECT 75.650 16.500 75.820 16.670 ;
        RECT 76.560 16.500 76.730 16.670 ;
        RECT 78.170 16.540 78.340 16.710 ;
        RECT 80.860 17.250 81.030 17.420 ;
        RECT 89.280 18.170 89.450 18.340 ;
        RECT 90.200 18.170 90.370 18.340 ;
        RECT 91.830 18.080 92.000 18.250 ;
        RECT 88.770 17.730 88.940 17.900 ;
        RECT 82.810 16.910 82.980 17.080 ;
        RECT 79.760 16.500 79.930 16.670 ;
        RECT 81.400 16.500 81.570 16.670 ;
        RECT 82.310 16.500 82.480 16.670 ;
        RECT 83.920 16.540 84.090 16.710 ;
        RECT 86.610 17.250 86.780 17.420 ;
        RECT 88.560 16.910 88.730 17.080 ;
        RECT 85.510 16.500 85.680 16.670 ;
        RECT 87.150 16.500 87.320 16.670 ;
        RECT 88.060 16.500 88.230 16.670 ;
        RECT 89.670 16.540 89.840 16.710 ;
        RECT 92.360 17.250 92.530 17.420 ;
        RECT 94.310 16.910 94.480 17.080 ;
        RECT 91.260 16.500 91.430 16.670 ;
        RECT 92.900 16.500 93.070 16.670 ;
        RECT 93.810 16.500 93.980 16.670 ;
        RECT 7.120 15.960 7.290 16.130 ;
        RECT 3.030 15.760 3.200 15.930 ;
        RECT 3.950 15.760 4.120 15.930 ;
        RECT 5.580 15.670 5.750 15.840 ;
        RECT 12.870 15.960 13.040 16.130 ;
        RECT 2.520 15.320 2.690 15.490 ;
        RECT 8.780 15.760 8.950 15.930 ;
        RECT 9.700 15.760 9.870 15.930 ;
        RECT 11.330 15.670 11.500 15.840 ;
        RECT 18.620 15.960 18.790 16.130 ;
        RECT 8.270 15.320 8.440 15.490 ;
        RECT 3.420 14.130 3.590 14.300 ;
        RECT 6.110 14.840 6.280 15.010 ;
        RECT 14.530 15.760 14.700 15.930 ;
        RECT 15.450 15.760 15.620 15.930 ;
        RECT 17.080 15.670 17.250 15.840 ;
        RECT 24.370 15.960 24.540 16.130 ;
        RECT 14.020 15.320 14.190 15.490 ;
        RECT 8.060 14.500 8.230 14.670 ;
        RECT 5.010 14.090 5.180 14.260 ;
        RECT 6.650 14.090 6.820 14.260 ;
        RECT 7.560 14.090 7.730 14.260 ;
        RECT 9.170 14.130 9.340 14.300 ;
        RECT 11.860 14.840 12.030 15.010 ;
        RECT 20.280 15.760 20.450 15.930 ;
        RECT 21.200 15.760 21.370 15.930 ;
        RECT 22.830 15.670 23.000 15.840 ;
        RECT 30.120 15.960 30.290 16.130 ;
        RECT 19.770 15.320 19.940 15.490 ;
        RECT 13.810 14.500 13.980 14.670 ;
        RECT 10.760 14.090 10.930 14.260 ;
        RECT 12.400 14.090 12.570 14.260 ;
        RECT 13.310 14.090 13.480 14.260 ;
        RECT 14.920 14.130 15.090 14.300 ;
        RECT 17.610 14.840 17.780 15.010 ;
        RECT 26.030 15.760 26.200 15.930 ;
        RECT 26.950 15.760 27.120 15.930 ;
        RECT 28.580 15.670 28.750 15.840 ;
        RECT 35.870 15.960 36.040 16.130 ;
        RECT 25.520 15.320 25.690 15.490 ;
        RECT 19.560 14.500 19.730 14.670 ;
        RECT 16.510 14.090 16.680 14.260 ;
        RECT 18.150 14.090 18.320 14.260 ;
        RECT 19.060 14.090 19.230 14.260 ;
        RECT 20.670 14.130 20.840 14.300 ;
        RECT 23.360 14.840 23.530 15.010 ;
        RECT 31.780 15.760 31.950 15.930 ;
        RECT 32.700 15.760 32.870 15.930 ;
        RECT 34.330 15.670 34.500 15.840 ;
        RECT 41.620 15.960 41.790 16.130 ;
        RECT 31.270 15.320 31.440 15.490 ;
        RECT 25.310 14.500 25.480 14.670 ;
        RECT 22.260 14.090 22.430 14.260 ;
        RECT 23.900 14.090 24.070 14.260 ;
        RECT 24.810 14.090 24.980 14.260 ;
        RECT 26.420 14.130 26.590 14.300 ;
        RECT 29.110 14.840 29.280 15.010 ;
        RECT 37.530 15.760 37.700 15.930 ;
        RECT 38.450 15.760 38.620 15.930 ;
        RECT 40.080 15.670 40.250 15.840 ;
        RECT 47.370 15.960 47.540 16.130 ;
        RECT 37.020 15.320 37.190 15.490 ;
        RECT 31.060 14.500 31.230 14.670 ;
        RECT 28.010 14.090 28.180 14.260 ;
        RECT 29.650 14.090 29.820 14.260 ;
        RECT 30.560 14.090 30.730 14.260 ;
        RECT 32.170 14.130 32.340 14.300 ;
        RECT 34.860 14.840 35.030 15.010 ;
        RECT 43.280 15.760 43.450 15.930 ;
        RECT 44.200 15.760 44.370 15.930 ;
        RECT 45.830 15.670 46.000 15.840 ;
        RECT 53.120 15.960 53.290 16.130 ;
        RECT 42.770 15.320 42.940 15.490 ;
        RECT 36.810 14.500 36.980 14.670 ;
        RECT 33.760 14.090 33.930 14.260 ;
        RECT 35.400 14.090 35.570 14.260 ;
        RECT 36.310 14.090 36.480 14.260 ;
        RECT 37.920 14.130 38.090 14.300 ;
        RECT 40.610 14.840 40.780 15.010 ;
        RECT 49.030 15.760 49.200 15.930 ;
        RECT 49.950 15.760 50.120 15.930 ;
        RECT 51.580 15.670 51.750 15.840 ;
        RECT 58.870 15.960 59.040 16.130 ;
        RECT 48.520 15.320 48.690 15.490 ;
        RECT 42.560 14.500 42.730 14.670 ;
        RECT 39.510 14.090 39.680 14.260 ;
        RECT 41.150 14.090 41.320 14.260 ;
        RECT 42.060 14.090 42.230 14.260 ;
        RECT 43.670 14.130 43.840 14.300 ;
        RECT 46.360 14.840 46.530 15.010 ;
        RECT 54.780 15.760 54.950 15.930 ;
        RECT 55.700 15.760 55.870 15.930 ;
        RECT 57.330 15.670 57.500 15.840 ;
        RECT 64.620 15.960 64.790 16.130 ;
        RECT 54.270 15.320 54.440 15.490 ;
        RECT 48.310 14.500 48.480 14.670 ;
        RECT 45.260 14.090 45.430 14.260 ;
        RECT 46.900 14.090 47.070 14.260 ;
        RECT 47.810 14.090 47.980 14.260 ;
        RECT 49.420 14.130 49.590 14.300 ;
        RECT 52.110 14.840 52.280 15.010 ;
        RECT 60.530 15.760 60.700 15.930 ;
        RECT 61.450 15.760 61.620 15.930 ;
        RECT 63.080 15.670 63.250 15.840 ;
        RECT 70.370 15.960 70.540 16.130 ;
        RECT 60.020 15.320 60.190 15.490 ;
        RECT 54.060 14.500 54.230 14.670 ;
        RECT 51.010 14.090 51.180 14.260 ;
        RECT 52.650 14.090 52.820 14.260 ;
        RECT 53.560 14.090 53.730 14.260 ;
        RECT 55.170 14.130 55.340 14.300 ;
        RECT 57.860 14.840 58.030 15.010 ;
        RECT 66.280 15.760 66.450 15.930 ;
        RECT 67.200 15.760 67.370 15.930 ;
        RECT 68.830 15.670 69.000 15.840 ;
        RECT 76.120 15.960 76.290 16.130 ;
        RECT 65.770 15.320 65.940 15.490 ;
        RECT 59.810 14.500 59.980 14.670 ;
        RECT 56.760 14.090 56.930 14.260 ;
        RECT 58.400 14.090 58.570 14.260 ;
        RECT 59.310 14.090 59.480 14.260 ;
        RECT 60.920 14.130 61.090 14.300 ;
        RECT 63.610 14.840 63.780 15.010 ;
        RECT 72.030 15.760 72.200 15.930 ;
        RECT 72.950 15.760 73.120 15.930 ;
        RECT 74.580 15.670 74.750 15.840 ;
        RECT 81.870 15.960 82.040 16.130 ;
        RECT 71.520 15.320 71.690 15.490 ;
        RECT 65.560 14.500 65.730 14.670 ;
        RECT 62.510 14.090 62.680 14.260 ;
        RECT 64.150 14.090 64.320 14.260 ;
        RECT 65.060 14.090 65.230 14.260 ;
        RECT 66.670 14.130 66.840 14.300 ;
        RECT 69.360 14.840 69.530 15.010 ;
        RECT 77.780 15.760 77.950 15.930 ;
        RECT 78.700 15.760 78.870 15.930 ;
        RECT 80.330 15.670 80.500 15.840 ;
        RECT 87.620 15.960 87.790 16.130 ;
        RECT 77.270 15.320 77.440 15.490 ;
        RECT 71.310 14.500 71.480 14.670 ;
        RECT 68.260 14.090 68.430 14.260 ;
        RECT 69.900 14.090 70.070 14.260 ;
        RECT 70.810 14.090 70.980 14.260 ;
        RECT 72.420 14.130 72.590 14.300 ;
        RECT 75.110 14.840 75.280 15.010 ;
        RECT 83.530 15.760 83.700 15.930 ;
        RECT 84.450 15.760 84.620 15.930 ;
        RECT 86.080 15.670 86.250 15.840 ;
        RECT 93.370 15.960 93.540 16.130 ;
        RECT 83.020 15.320 83.190 15.490 ;
        RECT 77.060 14.500 77.230 14.670 ;
        RECT 74.010 14.090 74.180 14.260 ;
        RECT 75.650 14.090 75.820 14.260 ;
        RECT 76.560 14.090 76.730 14.260 ;
        RECT 78.170 14.130 78.340 14.300 ;
        RECT 80.860 14.840 81.030 15.010 ;
        RECT 89.280 15.760 89.450 15.930 ;
        RECT 90.200 15.760 90.370 15.930 ;
        RECT 91.830 15.670 92.000 15.840 ;
        RECT 88.770 15.320 88.940 15.490 ;
        RECT 82.810 14.500 82.980 14.670 ;
        RECT 79.760 14.090 79.930 14.260 ;
        RECT 81.400 14.090 81.570 14.260 ;
        RECT 82.310 14.090 82.480 14.260 ;
        RECT 83.920 14.130 84.090 14.300 ;
        RECT 86.610 14.840 86.780 15.010 ;
        RECT 88.560 14.500 88.730 14.670 ;
        RECT 85.510 14.090 85.680 14.260 ;
        RECT 87.150 14.090 87.320 14.260 ;
        RECT 88.060 14.090 88.230 14.260 ;
        RECT 89.670 14.130 89.840 14.300 ;
        RECT 92.360 14.840 92.530 15.010 ;
        RECT 94.310 14.500 94.480 14.670 ;
        RECT 91.260 14.090 91.430 14.260 ;
        RECT 92.900 14.090 93.070 14.260 ;
        RECT 93.810 14.090 93.980 14.260 ;
        RECT 7.120 13.550 7.290 13.720 ;
        RECT 3.030 13.350 3.200 13.520 ;
        RECT 3.950 13.350 4.120 13.520 ;
        RECT 5.580 13.260 5.750 13.430 ;
        RECT 12.870 13.550 13.040 13.720 ;
        RECT 2.520 12.910 2.690 13.080 ;
        RECT 8.780 13.350 8.950 13.520 ;
        RECT 9.700 13.350 9.870 13.520 ;
        RECT 11.330 13.260 11.500 13.430 ;
        RECT 18.620 13.550 18.790 13.720 ;
        RECT 8.270 12.910 8.440 13.080 ;
        RECT 3.420 11.720 3.590 11.890 ;
        RECT 6.110 12.430 6.280 12.600 ;
        RECT 14.530 13.350 14.700 13.520 ;
        RECT 15.450 13.350 15.620 13.520 ;
        RECT 17.080 13.260 17.250 13.430 ;
        RECT 24.370 13.550 24.540 13.720 ;
        RECT 14.020 12.910 14.190 13.080 ;
        RECT 8.060 12.090 8.230 12.260 ;
        RECT 5.010 11.680 5.180 11.850 ;
        RECT 6.650 11.680 6.820 11.850 ;
        RECT 7.560 11.680 7.730 11.850 ;
        RECT 9.170 11.720 9.340 11.890 ;
        RECT 11.860 12.430 12.030 12.600 ;
        RECT 20.280 13.350 20.450 13.520 ;
        RECT 21.200 13.350 21.370 13.520 ;
        RECT 22.830 13.260 23.000 13.430 ;
        RECT 30.120 13.550 30.290 13.720 ;
        RECT 19.770 12.910 19.940 13.080 ;
        RECT 13.810 12.090 13.980 12.260 ;
        RECT 10.760 11.680 10.930 11.850 ;
        RECT 12.400 11.680 12.570 11.850 ;
        RECT 13.310 11.680 13.480 11.850 ;
        RECT 14.920 11.720 15.090 11.890 ;
        RECT 17.610 12.430 17.780 12.600 ;
        RECT 26.030 13.350 26.200 13.520 ;
        RECT 26.950 13.350 27.120 13.520 ;
        RECT 28.580 13.260 28.750 13.430 ;
        RECT 35.870 13.550 36.040 13.720 ;
        RECT 25.520 12.910 25.690 13.080 ;
        RECT 19.560 12.090 19.730 12.260 ;
        RECT 16.510 11.680 16.680 11.850 ;
        RECT 18.150 11.680 18.320 11.850 ;
        RECT 19.060 11.680 19.230 11.850 ;
        RECT 20.670 11.720 20.840 11.890 ;
        RECT 23.360 12.430 23.530 12.600 ;
        RECT 31.780 13.350 31.950 13.520 ;
        RECT 32.700 13.350 32.870 13.520 ;
        RECT 34.330 13.260 34.500 13.430 ;
        RECT 41.620 13.550 41.790 13.720 ;
        RECT 31.270 12.910 31.440 13.080 ;
        RECT 25.310 12.090 25.480 12.260 ;
        RECT 22.260 11.680 22.430 11.850 ;
        RECT 23.900 11.680 24.070 11.850 ;
        RECT 24.810 11.680 24.980 11.850 ;
        RECT 26.420 11.720 26.590 11.890 ;
        RECT 29.110 12.430 29.280 12.600 ;
        RECT 37.530 13.350 37.700 13.520 ;
        RECT 38.450 13.350 38.620 13.520 ;
        RECT 40.080 13.260 40.250 13.430 ;
        RECT 47.370 13.550 47.540 13.720 ;
        RECT 37.020 12.910 37.190 13.080 ;
        RECT 31.060 12.090 31.230 12.260 ;
        RECT 28.010 11.680 28.180 11.850 ;
        RECT 29.650 11.680 29.820 11.850 ;
        RECT 30.560 11.680 30.730 11.850 ;
        RECT 32.170 11.720 32.340 11.890 ;
        RECT 34.860 12.430 35.030 12.600 ;
        RECT 43.280 13.350 43.450 13.520 ;
        RECT 44.200 13.350 44.370 13.520 ;
        RECT 45.830 13.260 46.000 13.430 ;
        RECT 53.120 13.550 53.290 13.720 ;
        RECT 42.770 12.910 42.940 13.080 ;
        RECT 36.810 12.090 36.980 12.260 ;
        RECT 33.760 11.680 33.930 11.850 ;
        RECT 35.400 11.680 35.570 11.850 ;
        RECT 36.310 11.680 36.480 11.850 ;
        RECT 37.920 11.720 38.090 11.890 ;
        RECT 40.610 12.430 40.780 12.600 ;
        RECT 49.030 13.350 49.200 13.520 ;
        RECT 49.950 13.350 50.120 13.520 ;
        RECT 51.580 13.260 51.750 13.430 ;
        RECT 58.870 13.550 59.040 13.720 ;
        RECT 48.520 12.910 48.690 13.080 ;
        RECT 42.560 12.090 42.730 12.260 ;
        RECT 39.510 11.680 39.680 11.850 ;
        RECT 41.150 11.680 41.320 11.850 ;
        RECT 42.060 11.680 42.230 11.850 ;
        RECT 43.670 11.720 43.840 11.890 ;
        RECT 46.360 12.430 46.530 12.600 ;
        RECT 54.780 13.350 54.950 13.520 ;
        RECT 55.700 13.350 55.870 13.520 ;
        RECT 57.330 13.260 57.500 13.430 ;
        RECT 64.620 13.550 64.790 13.720 ;
        RECT 54.270 12.910 54.440 13.080 ;
        RECT 48.310 12.090 48.480 12.260 ;
        RECT 45.260 11.680 45.430 11.850 ;
        RECT 46.900 11.680 47.070 11.850 ;
        RECT 47.810 11.680 47.980 11.850 ;
        RECT 49.420 11.720 49.590 11.890 ;
        RECT 52.110 12.430 52.280 12.600 ;
        RECT 60.530 13.350 60.700 13.520 ;
        RECT 61.450 13.350 61.620 13.520 ;
        RECT 63.080 13.260 63.250 13.430 ;
        RECT 70.370 13.550 70.540 13.720 ;
        RECT 60.020 12.910 60.190 13.080 ;
        RECT 54.060 12.090 54.230 12.260 ;
        RECT 51.010 11.680 51.180 11.850 ;
        RECT 52.650 11.680 52.820 11.850 ;
        RECT 53.560 11.680 53.730 11.850 ;
        RECT 55.170 11.720 55.340 11.890 ;
        RECT 57.860 12.430 58.030 12.600 ;
        RECT 66.280 13.350 66.450 13.520 ;
        RECT 67.200 13.350 67.370 13.520 ;
        RECT 68.830 13.260 69.000 13.430 ;
        RECT 76.120 13.550 76.290 13.720 ;
        RECT 65.770 12.910 65.940 13.080 ;
        RECT 59.810 12.090 59.980 12.260 ;
        RECT 56.760 11.680 56.930 11.850 ;
        RECT 58.400 11.680 58.570 11.850 ;
        RECT 59.310 11.680 59.480 11.850 ;
        RECT 60.920 11.720 61.090 11.890 ;
        RECT 63.610 12.430 63.780 12.600 ;
        RECT 72.030 13.350 72.200 13.520 ;
        RECT 72.950 13.350 73.120 13.520 ;
        RECT 74.580 13.260 74.750 13.430 ;
        RECT 81.870 13.550 82.040 13.720 ;
        RECT 71.520 12.910 71.690 13.080 ;
        RECT 65.560 12.090 65.730 12.260 ;
        RECT 62.510 11.680 62.680 11.850 ;
        RECT 64.150 11.680 64.320 11.850 ;
        RECT 65.060 11.680 65.230 11.850 ;
        RECT 66.670 11.720 66.840 11.890 ;
        RECT 69.360 12.430 69.530 12.600 ;
        RECT 77.780 13.350 77.950 13.520 ;
        RECT 78.700 13.350 78.870 13.520 ;
        RECT 80.330 13.260 80.500 13.430 ;
        RECT 87.620 13.550 87.790 13.720 ;
        RECT 77.270 12.910 77.440 13.080 ;
        RECT 71.310 12.090 71.480 12.260 ;
        RECT 68.260 11.680 68.430 11.850 ;
        RECT 69.900 11.680 70.070 11.850 ;
        RECT 70.810 11.680 70.980 11.850 ;
        RECT 72.420 11.720 72.590 11.890 ;
        RECT 75.110 12.430 75.280 12.600 ;
        RECT 83.530 13.350 83.700 13.520 ;
        RECT 84.450 13.350 84.620 13.520 ;
        RECT 86.080 13.260 86.250 13.430 ;
        RECT 93.370 13.550 93.540 13.720 ;
        RECT 83.020 12.910 83.190 13.080 ;
        RECT 77.060 12.090 77.230 12.260 ;
        RECT 74.010 11.680 74.180 11.850 ;
        RECT 75.650 11.680 75.820 11.850 ;
        RECT 76.560 11.680 76.730 11.850 ;
        RECT 78.170 11.720 78.340 11.890 ;
        RECT 80.860 12.430 81.030 12.600 ;
        RECT 89.280 13.350 89.450 13.520 ;
        RECT 90.200 13.350 90.370 13.520 ;
        RECT 91.830 13.260 92.000 13.430 ;
        RECT 88.770 12.910 88.940 13.080 ;
        RECT 82.810 12.090 82.980 12.260 ;
        RECT 79.760 11.680 79.930 11.850 ;
        RECT 81.400 11.680 81.570 11.850 ;
        RECT 82.310 11.680 82.480 11.850 ;
        RECT 83.920 11.720 84.090 11.890 ;
        RECT 86.610 12.430 86.780 12.600 ;
        RECT 88.560 12.090 88.730 12.260 ;
        RECT 85.510 11.680 85.680 11.850 ;
        RECT 87.150 11.680 87.320 11.850 ;
        RECT 88.060 11.680 88.230 11.850 ;
        RECT 89.670 11.720 89.840 11.890 ;
        RECT 92.360 12.430 92.530 12.600 ;
        RECT 94.310 12.090 94.480 12.260 ;
        RECT 91.260 11.680 91.430 11.850 ;
        RECT 92.900 11.680 93.070 11.850 ;
        RECT 93.810 11.680 93.980 11.850 ;
        RECT 7.120 11.140 7.290 11.310 ;
        RECT 3.030 10.940 3.200 11.110 ;
        RECT 3.950 10.940 4.120 11.110 ;
        RECT 5.580 10.850 5.750 11.020 ;
        RECT 12.870 11.140 13.040 11.310 ;
        RECT 2.520 10.500 2.690 10.670 ;
        RECT 8.780 10.940 8.950 11.110 ;
        RECT 9.700 10.940 9.870 11.110 ;
        RECT 11.330 10.850 11.500 11.020 ;
        RECT 18.620 11.140 18.790 11.310 ;
        RECT 8.270 10.500 8.440 10.670 ;
        RECT 3.420 9.310 3.590 9.480 ;
        RECT 6.110 10.020 6.280 10.190 ;
        RECT 14.530 10.940 14.700 11.110 ;
        RECT 15.450 10.940 15.620 11.110 ;
        RECT 17.080 10.850 17.250 11.020 ;
        RECT 24.370 11.140 24.540 11.310 ;
        RECT 14.020 10.500 14.190 10.670 ;
        RECT 8.060 9.680 8.230 9.850 ;
        RECT 5.010 9.270 5.180 9.440 ;
        RECT 6.650 9.270 6.820 9.440 ;
        RECT 7.560 9.270 7.730 9.440 ;
        RECT 7.120 8.410 7.290 8.580 ;
        RECT 9.170 9.310 9.340 9.480 ;
        RECT 11.860 10.020 12.030 10.190 ;
        RECT 20.280 10.940 20.450 11.110 ;
        RECT 21.200 10.940 21.370 11.110 ;
        RECT 22.830 10.850 23.000 11.020 ;
        RECT 30.120 11.140 30.290 11.310 ;
        RECT 19.770 10.500 19.940 10.670 ;
        RECT 13.810 9.680 13.980 9.850 ;
        RECT 10.760 9.270 10.930 9.440 ;
        RECT 12.400 9.270 12.570 9.440 ;
        RECT 13.310 9.270 13.480 9.440 ;
        RECT 3.030 8.120 3.200 8.290 ;
        RECT 3.950 8.120 4.120 8.290 ;
        RECT 5.580 8.030 5.750 8.200 ;
        RECT 12.870 8.410 13.040 8.580 ;
        RECT 14.920 9.310 15.090 9.480 ;
        RECT 17.610 10.020 17.780 10.190 ;
        RECT 26.030 10.940 26.200 11.110 ;
        RECT 26.950 10.940 27.120 11.110 ;
        RECT 28.580 10.850 28.750 11.020 ;
        RECT 35.870 11.140 36.040 11.310 ;
        RECT 25.520 10.500 25.690 10.670 ;
        RECT 19.560 9.680 19.730 9.850 ;
        RECT 16.510 9.270 16.680 9.440 ;
        RECT 18.150 9.270 18.320 9.440 ;
        RECT 19.060 9.270 19.230 9.440 ;
        RECT 2.520 7.680 2.690 7.850 ;
        RECT 8.780 8.120 8.950 8.290 ;
        RECT 9.700 8.120 9.870 8.290 ;
        RECT 11.330 8.030 11.500 8.200 ;
        RECT 18.620 8.410 18.790 8.580 ;
        RECT 20.670 9.310 20.840 9.480 ;
        RECT 23.360 10.020 23.530 10.190 ;
        RECT 31.780 10.940 31.950 11.110 ;
        RECT 32.700 10.940 32.870 11.110 ;
        RECT 34.330 10.850 34.500 11.020 ;
        RECT 41.620 11.140 41.790 11.310 ;
        RECT 31.270 10.500 31.440 10.670 ;
        RECT 25.310 9.680 25.480 9.850 ;
        RECT 22.260 9.270 22.430 9.440 ;
        RECT 23.900 9.270 24.070 9.440 ;
        RECT 24.810 9.270 24.980 9.440 ;
        RECT 8.270 7.680 8.440 7.850 ;
        RECT 3.420 6.490 3.590 6.660 ;
        RECT 6.110 7.200 6.280 7.370 ;
        RECT 14.530 8.120 14.700 8.290 ;
        RECT 15.450 8.120 15.620 8.290 ;
        RECT 17.080 8.030 17.250 8.200 ;
        RECT 24.370 8.410 24.540 8.580 ;
        RECT 26.420 9.310 26.590 9.480 ;
        RECT 29.110 10.020 29.280 10.190 ;
        RECT 37.530 10.940 37.700 11.110 ;
        RECT 38.450 10.940 38.620 11.110 ;
        RECT 40.080 10.850 40.250 11.020 ;
        RECT 47.370 11.140 47.540 11.310 ;
        RECT 37.020 10.500 37.190 10.670 ;
        RECT 31.060 9.680 31.230 9.850 ;
        RECT 28.010 9.270 28.180 9.440 ;
        RECT 29.650 9.270 29.820 9.440 ;
        RECT 30.560 9.270 30.730 9.440 ;
        RECT 14.020 7.680 14.190 7.850 ;
        RECT 8.060 6.860 8.230 7.030 ;
        RECT 5.010 6.450 5.180 6.620 ;
        RECT 6.650 6.450 6.820 6.620 ;
        RECT 7.560 6.450 7.730 6.620 ;
        RECT 9.170 6.490 9.340 6.660 ;
        RECT 11.860 7.200 12.030 7.370 ;
        RECT 20.280 8.120 20.450 8.290 ;
        RECT 21.200 8.120 21.370 8.290 ;
        RECT 22.830 8.030 23.000 8.200 ;
        RECT 30.120 8.410 30.290 8.580 ;
        RECT 32.170 9.310 32.340 9.480 ;
        RECT 34.860 10.020 35.030 10.190 ;
        RECT 43.280 10.940 43.450 11.110 ;
        RECT 44.200 10.940 44.370 11.110 ;
        RECT 45.830 10.850 46.000 11.020 ;
        RECT 53.120 11.140 53.290 11.310 ;
        RECT 42.770 10.500 42.940 10.670 ;
        RECT 36.810 9.680 36.980 9.850 ;
        RECT 33.760 9.270 33.930 9.440 ;
        RECT 35.400 9.270 35.570 9.440 ;
        RECT 36.310 9.270 36.480 9.440 ;
        RECT 19.770 7.680 19.940 7.850 ;
        RECT 13.810 6.860 13.980 7.030 ;
        RECT 10.760 6.450 10.930 6.620 ;
        RECT 12.400 6.450 12.570 6.620 ;
        RECT 13.310 6.450 13.480 6.620 ;
        RECT 14.920 6.490 15.090 6.660 ;
        RECT 17.610 7.200 17.780 7.370 ;
        RECT 26.030 8.120 26.200 8.290 ;
        RECT 26.950 8.120 27.120 8.290 ;
        RECT 28.580 8.030 28.750 8.200 ;
        RECT 35.870 8.410 36.040 8.580 ;
        RECT 37.920 9.310 38.090 9.480 ;
        RECT 40.610 10.020 40.780 10.190 ;
        RECT 49.030 10.940 49.200 11.110 ;
        RECT 49.950 10.940 50.120 11.110 ;
        RECT 51.580 10.850 51.750 11.020 ;
        RECT 58.870 11.140 59.040 11.310 ;
        RECT 48.520 10.500 48.690 10.670 ;
        RECT 42.560 9.680 42.730 9.850 ;
        RECT 39.510 9.270 39.680 9.440 ;
        RECT 41.150 9.270 41.320 9.440 ;
        RECT 42.060 9.270 42.230 9.440 ;
        RECT 25.520 7.680 25.690 7.850 ;
        RECT 19.560 6.860 19.730 7.030 ;
        RECT 16.510 6.450 16.680 6.620 ;
        RECT 18.150 6.450 18.320 6.620 ;
        RECT 19.060 6.450 19.230 6.620 ;
        RECT 20.670 6.490 20.840 6.660 ;
        RECT 23.360 7.200 23.530 7.370 ;
        RECT 31.780 8.120 31.950 8.290 ;
        RECT 32.700 8.120 32.870 8.290 ;
        RECT 34.330 8.030 34.500 8.200 ;
        RECT 41.620 8.410 41.790 8.580 ;
        RECT 43.670 9.310 43.840 9.480 ;
        RECT 46.360 10.020 46.530 10.190 ;
        RECT 54.780 10.940 54.950 11.110 ;
        RECT 55.700 10.940 55.870 11.110 ;
        RECT 57.330 10.850 57.500 11.020 ;
        RECT 64.620 11.140 64.790 11.310 ;
        RECT 54.270 10.500 54.440 10.670 ;
        RECT 48.310 9.680 48.480 9.850 ;
        RECT 45.260 9.270 45.430 9.440 ;
        RECT 46.900 9.270 47.070 9.440 ;
        RECT 47.810 9.270 47.980 9.440 ;
        RECT 31.270 7.680 31.440 7.850 ;
        RECT 25.310 6.860 25.480 7.030 ;
        RECT 22.260 6.450 22.430 6.620 ;
        RECT 23.900 6.450 24.070 6.620 ;
        RECT 24.810 6.450 24.980 6.620 ;
        RECT 26.420 6.490 26.590 6.660 ;
        RECT 29.110 7.200 29.280 7.370 ;
        RECT 37.530 8.120 37.700 8.290 ;
        RECT 38.450 8.120 38.620 8.290 ;
        RECT 40.080 8.030 40.250 8.200 ;
        RECT 47.370 8.410 47.540 8.580 ;
        RECT 49.420 9.310 49.590 9.480 ;
        RECT 52.110 10.020 52.280 10.190 ;
        RECT 60.530 10.940 60.700 11.110 ;
        RECT 61.450 10.940 61.620 11.110 ;
        RECT 63.080 10.850 63.250 11.020 ;
        RECT 70.370 11.140 70.540 11.310 ;
        RECT 60.020 10.500 60.190 10.670 ;
        RECT 54.060 9.680 54.230 9.850 ;
        RECT 51.010 9.270 51.180 9.440 ;
        RECT 52.650 9.270 52.820 9.440 ;
        RECT 53.560 9.270 53.730 9.440 ;
        RECT 37.020 7.680 37.190 7.850 ;
        RECT 31.060 6.860 31.230 7.030 ;
        RECT 28.010 6.450 28.180 6.620 ;
        RECT 29.650 6.450 29.820 6.620 ;
        RECT 30.560 6.450 30.730 6.620 ;
        RECT 32.170 6.490 32.340 6.660 ;
        RECT 34.860 7.200 35.030 7.370 ;
        RECT 43.280 8.120 43.450 8.290 ;
        RECT 44.200 8.120 44.370 8.290 ;
        RECT 45.830 8.030 46.000 8.200 ;
        RECT 53.120 8.410 53.290 8.580 ;
        RECT 55.170 9.310 55.340 9.480 ;
        RECT 57.860 10.020 58.030 10.190 ;
        RECT 66.280 10.940 66.450 11.110 ;
        RECT 67.200 10.940 67.370 11.110 ;
        RECT 68.830 10.850 69.000 11.020 ;
        RECT 76.120 11.140 76.290 11.310 ;
        RECT 65.770 10.500 65.940 10.670 ;
        RECT 59.810 9.680 59.980 9.850 ;
        RECT 56.760 9.270 56.930 9.440 ;
        RECT 58.400 9.270 58.570 9.440 ;
        RECT 59.310 9.270 59.480 9.440 ;
        RECT 42.770 7.680 42.940 7.850 ;
        RECT 36.810 6.860 36.980 7.030 ;
        RECT 33.760 6.450 33.930 6.620 ;
        RECT 35.400 6.450 35.570 6.620 ;
        RECT 36.310 6.450 36.480 6.620 ;
        RECT 37.920 6.490 38.090 6.660 ;
        RECT 40.610 7.200 40.780 7.370 ;
        RECT 49.030 8.120 49.200 8.290 ;
        RECT 49.950 8.120 50.120 8.290 ;
        RECT 51.580 8.030 51.750 8.200 ;
        RECT 58.870 8.410 59.040 8.580 ;
        RECT 60.920 9.310 61.090 9.480 ;
        RECT 63.610 10.020 63.780 10.190 ;
        RECT 72.030 10.940 72.200 11.110 ;
        RECT 72.950 10.940 73.120 11.110 ;
        RECT 74.580 10.850 74.750 11.020 ;
        RECT 81.870 11.140 82.040 11.310 ;
        RECT 71.520 10.500 71.690 10.670 ;
        RECT 65.560 9.680 65.730 9.850 ;
        RECT 62.510 9.270 62.680 9.440 ;
        RECT 64.150 9.270 64.320 9.440 ;
        RECT 65.060 9.270 65.230 9.440 ;
        RECT 48.520 7.680 48.690 7.850 ;
        RECT 42.560 6.860 42.730 7.030 ;
        RECT 39.510 6.450 39.680 6.620 ;
        RECT 41.150 6.450 41.320 6.620 ;
        RECT 42.060 6.450 42.230 6.620 ;
        RECT 43.670 6.490 43.840 6.660 ;
        RECT 46.360 7.200 46.530 7.370 ;
        RECT 54.780 8.120 54.950 8.290 ;
        RECT 55.700 8.120 55.870 8.290 ;
        RECT 57.330 8.030 57.500 8.200 ;
        RECT 64.620 8.410 64.790 8.580 ;
        RECT 66.670 9.310 66.840 9.480 ;
        RECT 69.360 10.020 69.530 10.190 ;
        RECT 77.780 10.940 77.950 11.110 ;
        RECT 78.700 10.940 78.870 11.110 ;
        RECT 80.330 10.850 80.500 11.020 ;
        RECT 87.620 11.140 87.790 11.310 ;
        RECT 77.270 10.500 77.440 10.670 ;
        RECT 71.310 9.680 71.480 9.850 ;
        RECT 68.260 9.270 68.430 9.440 ;
        RECT 69.900 9.270 70.070 9.440 ;
        RECT 70.810 9.270 70.980 9.440 ;
        RECT 54.270 7.680 54.440 7.850 ;
        RECT 48.310 6.860 48.480 7.030 ;
        RECT 45.260 6.450 45.430 6.620 ;
        RECT 46.900 6.450 47.070 6.620 ;
        RECT 47.810 6.450 47.980 6.620 ;
        RECT 49.420 6.490 49.590 6.660 ;
        RECT 52.110 7.200 52.280 7.370 ;
        RECT 60.530 8.120 60.700 8.290 ;
        RECT 61.450 8.120 61.620 8.290 ;
        RECT 63.080 8.030 63.250 8.200 ;
        RECT 70.370 8.410 70.540 8.580 ;
        RECT 72.420 9.310 72.590 9.480 ;
        RECT 75.110 10.020 75.280 10.190 ;
        RECT 83.530 10.940 83.700 11.110 ;
        RECT 84.450 10.940 84.620 11.110 ;
        RECT 86.080 10.850 86.250 11.020 ;
        RECT 93.370 11.140 93.540 11.310 ;
        RECT 83.020 10.500 83.190 10.670 ;
        RECT 77.060 9.680 77.230 9.850 ;
        RECT 74.010 9.270 74.180 9.440 ;
        RECT 75.650 9.270 75.820 9.440 ;
        RECT 76.560 9.270 76.730 9.440 ;
        RECT 60.020 7.680 60.190 7.850 ;
        RECT 54.060 6.860 54.230 7.030 ;
        RECT 51.010 6.450 51.180 6.620 ;
        RECT 52.650 6.450 52.820 6.620 ;
        RECT 53.560 6.450 53.730 6.620 ;
        RECT 55.170 6.490 55.340 6.660 ;
        RECT 57.860 7.200 58.030 7.370 ;
        RECT 66.280 8.120 66.450 8.290 ;
        RECT 67.200 8.120 67.370 8.290 ;
        RECT 68.830 8.030 69.000 8.200 ;
        RECT 76.120 8.410 76.290 8.580 ;
        RECT 78.170 9.310 78.340 9.480 ;
        RECT 80.860 10.020 81.030 10.190 ;
        RECT 89.280 10.940 89.450 11.110 ;
        RECT 90.200 10.940 90.370 11.110 ;
        RECT 91.830 10.850 92.000 11.020 ;
        RECT 88.770 10.500 88.940 10.670 ;
        RECT 82.810 9.680 82.980 9.850 ;
        RECT 79.760 9.270 79.930 9.440 ;
        RECT 81.400 9.270 81.570 9.440 ;
        RECT 82.310 9.270 82.480 9.440 ;
        RECT 65.770 7.680 65.940 7.850 ;
        RECT 59.810 6.860 59.980 7.030 ;
        RECT 56.760 6.450 56.930 6.620 ;
        RECT 58.400 6.450 58.570 6.620 ;
        RECT 59.310 6.450 59.480 6.620 ;
        RECT 60.920 6.490 61.090 6.660 ;
        RECT 63.610 7.200 63.780 7.370 ;
        RECT 72.030 8.120 72.200 8.290 ;
        RECT 72.950 8.120 73.120 8.290 ;
        RECT 74.580 8.030 74.750 8.200 ;
        RECT 81.870 8.410 82.040 8.580 ;
        RECT 83.920 9.310 84.090 9.480 ;
        RECT 86.610 10.020 86.780 10.190 ;
        RECT 88.560 9.680 88.730 9.850 ;
        RECT 85.510 9.270 85.680 9.440 ;
        RECT 87.150 9.270 87.320 9.440 ;
        RECT 88.060 9.270 88.230 9.440 ;
        RECT 71.520 7.680 71.690 7.850 ;
        RECT 65.560 6.860 65.730 7.030 ;
        RECT 62.510 6.450 62.680 6.620 ;
        RECT 64.150 6.450 64.320 6.620 ;
        RECT 65.060 6.450 65.230 6.620 ;
        RECT 66.670 6.490 66.840 6.660 ;
        RECT 69.360 7.200 69.530 7.370 ;
        RECT 77.780 8.120 77.950 8.290 ;
        RECT 78.700 8.120 78.870 8.290 ;
        RECT 80.330 8.030 80.500 8.200 ;
        RECT 87.620 8.410 87.790 8.580 ;
        RECT 89.670 9.310 89.840 9.480 ;
        RECT 92.360 10.020 92.530 10.190 ;
        RECT 94.310 9.680 94.480 9.850 ;
        RECT 91.260 9.270 91.430 9.440 ;
        RECT 92.900 9.270 93.070 9.440 ;
        RECT 93.810 9.270 93.980 9.440 ;
        RECT 77.270 7.680 77.440 7.850 ;
        RECT 71.310 6.860 71.480 7.030 ;
        RECT 68.260 6.450 68.430 6.620 ;
        RECT 69.900 6.450 70.070 6.620 ;
        RECT 70.810 6.450 70.980 6.620 ;
        RECT 72.420 6.490 72.590 6.660 ;
        RECT 75.110 7.200 75.280 7.370 ;
        RECT 83.530 8.120 83.700 8.290 ;
        RECT 84.450 8.120 84.620 8.290 ;
        RECT 86.080 8.030 86.250 8.200 ;
        RECT 83.020 7.680 83.190 7.850 ;
        RECT 77.060 6.860 77.230 7.030 ;
        RECT 74.010 6.450 74.180 6.620 ;
        RECT 75.650 6.450 75.820 6.620 ;
        RECT 76.560 6.450 76.730 6.620 ;
        RECT 78.170 6.490 78.340 6.660 ;
        RECT 80.860 7.200 81.030 7.370 ;
        RECT 89.280 8.120 89.450 8.290 ;
        RECT 90.200 8.120 90.370 8.290 ;
        RECT 91.830 8.030 92.000 8.200 ;
        RECT 88.770 7.680 88.940 7.850 ;
        RECT 82.810 6.860 82.980 7.030 ;
        RECT 79.760 6.450 79.930 6.620 ;
        RECT 81.400 6.450 81.570 6.620 ;
        RECT 82.310 6.450 82.480 6.620 ;
        RECT 83.920 6.490 84.090 6.660 ;
        RECT 86.610 7.200 86.780 7.370 ;
        RECT 88.560 6.860 88.730 7.030 ;
        RECT 85.510 6.450 85.680 6.620 ;
        RECT 87.150 6.450 87.320 6.620 ;
        RECT 88.060 6.450 88.230 6.620 ;
        RECT 89.670 6.490 89.840 6.660 ;
        RECT 92.360 7.200 92.530 7.370 ;
        RECT 94.310 6.860 94.480 7.030 ;
        RECT 91.260 6.450 91.430 6.620 ;
        RECT 92.900 6.450 93.070 6.620 ;
        RECT 93.810 6.450 93.980 6.620 ;
        RECT 7.120 5.910 7.290 6.080 ;
        RECT 3.030 5.710 3.200 5.880 ;
        RECT 3.950 5.710 4.120 5.880 ;
        RECT 5.580 5.620 5.750 5.790 ;
        RECT 12.870 5.910 13.040 6.080 ;
        RECT 2.520 5.270 2.690 5.440 ;
        RECT 8.780 5.710 8.950 5.880 ;
        RECT 9.700 5.710 9.870 5.880 ;
        RECT 11.330 5.620 11.500 5.790 ;
        RECT 18.620 5.910 18.790 6.080 ;
        RECT 8.270 5.270 8.440 5.440 ;
        RECT 3.420 4.080 3.590 4.250 ;
        RECT 6.110 4.790 6.280 4.960 ;
        RECT 14.530 5.710 14.700 5.880 ;
        RECT 15.450 5.710 15.620 5.880 ;
        RECT 17.080 5.620 17.250 5.790 ;
        RECT 24.370 5.910 24.540 6.080 ;
        RECT 14.020 5.270 14.190 5.440 ;
        RECT 8.060 4.450 8.230 4.620 ;
        RECT 5.010 4.040 5.180 4.210 ;
        RECT 6.650 4.040 6.820 4.210 ;
        RECT 7.560 4.040 7.730 4.210 ;
        RECT 9.170 4.080 9.340 4.250 ;
        RECT 11.860 4.790 12.030 4.960 ;
        RECT 20.280 5.710 20.450 5.880 ;
        RECT 21.200 5.710 21.370 5.880 ;
        RECT 22.830 5.620 23.000 5.790 ;
        RECT 30.120 5.910 30.290 6.080 ;
        RECT 19.770 5.270 19.940 5.440 ;
        RECT 13.810 4.450 13.980 4.620 ;
        RECT 10.760 4.040 10.930 4.210 ;
        RECT 12.400 4.040 12.570 4.210 ;
        RECT 13.310 4.040 13.480 4.210 ;
        RECT 14.920 4.080 15.090 4.250 ;
        RECT 17.610 4.790 17.780 4.960 ;
        RECT 26.030 5.710 26.200 5.880 ;
        RECT 26.950 5.710 27.120 5.880 ;
        RECT 28.580 5.620 28.750 5.790 ;
        RECT 35.870 5.910 36.040 6.080 ;
        RECT 25.520 5.270 25.690 5.440 ;
        RECT 19.560 4.450 19.730 4.620 ;
        RECT 16.510 4.040 16.680 4.210 ;
        RECT 18.150 4.040 18.320 4.210 ;
        RECT 19.060 4.040 19.230 4.210 ;
        RECT 20.670 4.080 20.840 4.250 ;
        RECT 23.360 4.790 23.530 4.960 ;
        RECT 31.780 5.710 31.950 5.880 ;
        RECT 32.700 5.710 32.870 5.880 ;
        RECT 34.330 5.620 34.500 5.790 ;
        RECT 41.620 5.910 41.790 6.080 ;
        RECT 31.270 5.270 31.440 5.440 ;
        RECT 25.310 4.450 25.480 4.620 ;
        RECT 22.260 4.040 22.430 4.210 ;
        RECT 23.900 4.040 24.070 4.210 ;
        RECT 24.810 4.040 24.980 4.210 ;
        RECT 26.420 4.080 26.590 4.250 ;
        RECT 29.110 4.790 29.280 4.960 ;
        RECT 37.530 5.710 37.700 5.880 ;
        RECT 38.450 5.710 38.620 5.880 ;
        RECT 40.080 5.620 40.250 5.790 ;
        RECT 47.370 5.910 47.540 6.080 ;
        RECT 37.020 5.270 37.190 5.440 ;
        RECT 31.060 4.450 31.230 4.620 ;
        RECT 28.010 4.040 28.180 4.210 ;
        RECT 29.650 4.040 29.820 4.210 ;
        RECT 30.560 4.040 30.730 4.210 ;
        RECT 32.170 4.080 32.340 4.250 ;
        RECT 34.860 4.790 35.030 4.960 ;
        RECT 43.280 5.710 43.450 5.880 ;
        RECT 44.200 5.710 44.370 5.880 ;
        RECT 45.830 5.620 46.000 5.790 ;
        RECT 53.120 5.910 53.290 6.080 ;
        RECT 42.770 5.270 42.940 5.440 ;
        RECT 36.810 4.450 36.980 4.620 ;
        RECT 33.760 4.040 33.930 4.210 ;
        RECT 35.400 4.040 35.570 4.210 ;
        RECT 36.310 4.040 36.480 4.210 ;
        RECT 37.920 4.080 38.090 4.250 ;
        RECT 40.610 4.790 40.780 4.960 ;
        RECT 49.030 5.710 49.200 5.880 ;
        RECT 49.950 5.710 50.120 5.880 ;
        RECT 51.580 5.620 51.750 5.790 ;
        RECT 58.870 5.910 59.040 6.080 ;
        RECT 48.520 5.270 48.690 5.440 ;
        RECT 42.560 4.450 42.730 4.620 ;
        RECT 39.510 4.040 39.680 4.210 ;
        RECT 41.150 4.040 41.320 4.210 ;
        RECT 42.060 4.040 42.230 4.210 ;
        RECT 43.670 4.080 43.840 4.250 ;
        RECT 46.360 4.790 46.530 4.960 ;
        RECT 54.780 5.710 54.950 5.880 ;
        RECT 55.700 5.710 55.870 5.880 ;
        RECT 57.330 5.620 57.500 5.790 ;
        RECT 64.620 5.910 64.790 6.080 ;
        RECT 54.270 5.270 54.440 5.440 ;
        RECT 48.310 4.450 48.480 4.620 ;
        RECT 45.260 4.040 45.430 4.210 ;
        RECT 46.900 4.040 47.070 4.210 ;
        RECT 47.810 4.040 47.980 4.210 ;
        RECT 49.420 4.080 49.590 4.250 ;
        RECT 52.110 4.790 52.280 4.960 ;
        RECT 60.530 5.710 60.700 5.880 ;
        RECT 61.450 5.710 61.620 5.880 ;
        RECT 63.080 5.620 63.250 5.790 ;
        RECT 70.370 5.910 70.540 6.080 ;
        RECT 60.020 5.270 60.190 5.440 ;
        RECT 54.060 4.450 54.230 4.620 ;
        RECT 51.010 4.040 51.180 4.210 ;
        RECT 52.650 4.040 52.820 4.210 ;
        RECT 53.560 4.040 53.730 4.210 ;
        RECT 55.170 4.080 55.340 4.250 ;
        RECT 57.860 4.790 58.030 4.960 ;
        RECT 66.280 5.710 66.450 5.880 ;
        RECT 67.200 5.710 67.370 5.880 ;
        RECT 68.830 5.620 69.000 5.790 ;
        RECT 76.120 5.910 76.290 6.080 ;
        RECT 65.770 5.270 65.940 5.440 ;
        RECT 59.810 4.450 59.980 4.620 ;
        RECT 56.760 4.040 56.930 4.210 ;
        RECT 58.400 4.040 58.570 4.210 ;
        RECT 59.310 4.040 59.480 4.210 ;
        RECT 60.920 4.080 61.090 4.250 ;
        RECT 63.610 4.790 63.780 4.960 ;
        RECT 72.030 5.710 72.200 5.880 ;
        RECT 72.950 5.710 73.120 5.880 ;
        RECT 74.580 5.620 74.750 5.790 ;
        RECT 81.870 5.910 82.040 6.080 ;
        RECT 71.520 5.270 71.690 5.440 ;
        RECT 65.560 4.450 65.730 4.620 ;
        RECT 62.510 4.040 62.680 4.210 ;
        RECT 64.150 4.040 64.320 4.210 ;
        RECT 65.060 4.040 65.230 4.210 ;
        RECT 66.670 4.080 66.840 4.250 ;
        RECT 69.360 4.790 69.530 4.960 ;
        RECT 77.780 5.710 77.950 5.880 ;
        RECT 78.700 5.710 78.870 5.880 ;
        RECT 80.330 5.620 80.500 5.790 ;
        RECT 87.620 5.910 87.790 6.080 ;
        RECT 77.270 5.270 77.440 5.440 ;
        RECT 71.310 4.450 71.480 4.620 ;
        RECT 68.260 4.040 68.430 4.210 ;
        RECT 69.900 4.040 70.070 4.210 ;
        RECT 70.810 4.040 70.980 4.210 ;
        RECT 72.420 4.080 72.590 4.250 ;
        RECT 75.110 4.790 75.280 4.960 ;
        RECT 83.530 5.710 83.700 5.880 ;
        RECT 84.450 5.710 84.620 5.880 ;
        RECT 86.080 5.620 86.250 5.790 ;
        RECT 93.370 5.910 93.540 6.080 ;
        RECT 83.020 5.270 83.190 5.440 ;
        RECT 77.060 4.450 77.230 4.620 ;
        RECT 74.010 4.040 74.180 4.210 ;
        RECT 75.650 4.040 75.820 4.210 ;
        RECT 76.560 4.040 76.730 4.210 ;
        RECT 78.170 4.080 78.340 4.250 ;
        RECT 80.860 4.790 81.030 4.960 ;
        RECT 89.280 5.710 89.450 5.880 ;
        RECT 90.200 5.710 90.370 5.880 ;
        RECT 91.830 5.620 92.000 5.790 ;
        RECT 88.770 5.270 88.940 5.440 ;
        RECT 82.810 4.450 82.980 4.620 ;
        RECT 79.760 4.040 79.930 4.210 ;
        RECT 81.400 4.040 81.570 4.210 ;
        RECT 82.310 4.040 82.480 4.210 ;
        RECT 83.920 4.080 84.090 4.250 ;
        RECT 86.610 4.790 86.780 4.960 ;
        RECT 88.560 4.450 88.730 4.620 ;
        RECT 85.510 4.040 85.680 4.210 ;
        RECT 87.150 4.040 87.320 4.210 ;
        RECT 88.060 4.040 88.230 4.210 ;
        RECT 89.670 4.080 89.840 4.250 ;
        RECT 92.360 4.790 92.530 4.960 ;
        RECT 94.310 4.450 94.480 4.620 ;
        RECT 91.260 4.040 91.430 4.210 ;
        RECT 92.900 4.040 93.070 4.210 ;
        RECT 93.810 4.040 93.980 4.210 ;
        RECT 7.120 3.500 7.290 3.670 ;
        RECT 3.030 3.300 3.200 3.470 ;
        RECT 3.950 3.300 4.120 3.470 ;
        RECT 5.580 3.210 5.750 3.380 ;
        RECT 12.870 3.500 13.040 3.670 ;
        RECT 2.520 2.860 2.690 3.030 ;
        RECT 8.780 3.300 8.950 3.470 ;
        RECT 9.700 3.300 9.870 3.470 ;
        RECT 11.330 3.210 11.500 3.380 ;
        RECT 18.620 3.500 18.790 3.670 ;
        RECT 8.270 2.860 8.440 3.030 ;
        RECT 3.420 1.670 3.590 1.840 ;
        RECT 6.110 2.380 6.280 2.550 ;
        RECT 14.530 3.300 14.700 3.470 ;
        RECT 15.450 3.300 15.620 3.470 ;
        RECT 17.080 3.210 17.250 3.380 ;
        RECT 24.370 3.500 24.540 3.670 ;
        RECT 14.020 2.860 14.190 3.030 ;
        RECT 8.060 2.040 8.230 2.210 ;
        RECT 5.010 1.630 5.180 1.800 ;
        RECT 6.650 1.630 6.820 1.800 ;
        RECT 7.560 1.630 7.730 1.800 ;
        RECT 9.170 1.670 9.340 1.840 ;
        RECT 11.860 2.380 12.030 2.550 ;
        RECT 20.280 3.300 20.450 3.470 ;
        RECT 21.200 3.300 21.370 3.470 ;
        RECT 22.830 3.210 23.000 3.380 ;
        RECT 30.120 3.500 30.290 3.670 ;
        RECT 19.770 2.860 19.940 3.030 ;
        RECT 13.810 2.040 13.980 2.210 ;
        RECT 10.760 1.630 10.930 1.800 ;
        RECT 12.400 1.630 12.570 1.800 ;
        RECT 13.310 1.630 13.480 1.800 ;
        RECT 14.920 1.670 15.090 1.840 ;
        RECT 17.610 2.380 17.780 2.550 ;
        RECT 26.030 3.300 26.200 3.470 ;
        RECT 26.950 3.300 27.120 3.470 ;
        RECT 28.580 3.210 28.750 3.380 ;
        RECT 35.870 3.500 36.040 3.670 ;
        RECT 25.520 2.860 25.690 3.030 ;
        RECT 19.560 2.040 19.730 2.210 ;
        RECT 16.510 1.630 16.680 1.800 ;
        RECT 18.150 1.630 18.320 1.800 ;
        RECT 19.060 1.630 19.230 1.800 ;
        RECT 20.670 1.670 20.840 1.840 ;
        RECT 23.360 2.380 23.530 2.550 ;
        RECT 31.780 3.300 31.950 3.470 ;
        RECT 32.700 3.300 32.870 3.470 ;
        RECT 34.330 3.210 34.500 3.380 ;
        RECT 41.620 3.500 41.790 3.670 ;
        RECT 31.270 2.860 31.440 3.030 ;
        RECT 25.310 2.040 25.480 2.210 ;
        RECT 22.260 1.630 22.430 1.800 ;
        RECT 23.900 1.630 24.070 1.800 ;
        RECT 24.810 1.630 24.980 1.800 ;
        RECT 26.420 1.670 26.590 1.840 ;
        RECT 29.110 2.380 29.280 2.550 ;
        RECT 37.530 3.300 37.700 3.470 ;
        RECT 38.450 3.300 38.620 3.470 ;
        RECT 40.080 3.210 40.250 3.380 ;
        RECT 47.370 3.500 47.540 3.670 ;
        RECT 37.020 2.860 37.190 3.030 ;
        RECT 31.060 2.040 31.230 2.210 ;
        RECT 28.010 1.630 28.180 1.800 ;
        RECT 29.650 1.630 29.820 1.800 ;
        RECT 30.560 1.630 30.730 1.800 ;
        RECT 32.170 1.670 32.340 1.840 ;
        RECT 34.860 2.380 35.030 2.550 ;
        RECT 43.280 3.300 43.450 3.470 ;
        RECT 44.200 3.300 44.370 3.470 ;
        RECT 45.830 3.210 46.000 3.380 ;
        RECT 53.120 3.500 53.290 3.670 ;
        RECT 42.770 2.860 42.940 3.030 ;
        RECT 36.810 2.040 36.980 2.210 ;
        RECT 33.760 1.630 33.930 1.800 ;
        RECT 35.400 1.630 35.570 1.800 ;
        RECT 36.310 1.630 36.480 1.800 ;
        RECT 37.920 1.670 38.090 1.840 ;
        RECT 40.610 2.380 40.780 2.550 ;
        RECT 49.030 3.300 49.200 3.470 ;
        RECT 49.950 3.300 50.120 3.470 ;
        RECT 51.580 3.210 51.750 3.380 ;
        RECT 58.870 3.500 59.040 3.670 ;
        RECT 48.520 2.860 48.690 3.030 ;
        RECT 42.560 2.040 42.730 2.210 ;
        RECT 39.510 1.630 39.680 1.800 ;
        RECT 41.150 1.630 41.320 1.800 ;
        RECT 42.060 1.630 42.230 1.800 ;
        RECT 43.670 1.670 43.840 1.840 ;
        RECT 46.360 2.380 46.530 2.550 ;
        RECT 54.780 3.300 54.950 3.470 ;
        RECT 55.700 3.300 55.870 3.470 ;
        RECT 57.330 3.210 57.500 3.380 ;
        RECT 64.620 3.500 64.790 3.670 ;
        RECT 54.270 2.860 54.440 3.030 ;
        RECT 48.310 2.040 48.480 2.210 ;
        RECT 45.260 1.630 45.430 1.800 ;
        RECT 46.900 1.630 47.070 1.800 ;
        RECT 47.810 1.630 47.980 1.800 ;
        RECT 49.420 1.670 49.590 1.840 ;
        RECT 52.110 2.380 52.280 2.550 ;
        RECT 60.530 3.300 60.700 3.470 ;
        RECT 61.450 3.300 61.620 3.470 ;
        RECT 63.080 3.210 63.250 3.380 ;
        RECT 70.370 3.500 70.540 3.670 ;
        RECT 60.020 2.860 60.190 3.030 ;
        RECT 54.060 2.040 54.230 2.210 ;
        RECT 51.010 1.630 51.180 1.800 ;
        RECT 52.650 1.630 52.820 1.800 ;
        RECT 53.560 1.630 53.730 1.800 ;
        RECT 55.170 1.670 55.340 1.840 ;
        RECT 57.860 2.380 58.030 2.550 ;
        RECT 66.280 3.300 66.450 3.470 ;
        RECT 67.200 3.300 67.370 3.470 ;
        RECT 68.830 3.210 69.000 3.380 ;
        RECT 76.120 3.500 76.290 3.670 ;
        RECT 65.770 2.860 65.940 3.030 ;
        RECT 59.810 2.040 59.980 2.210 ;
        RECT 56.760 1.630 56.930 1.800 ;
        RECT 58.400 1.630 58.570 1.800 ;
        RECT 59.310 1.630 59.480 1.800 ;
        RECT 60.920 1.670 61.090 1.840 ;
        RECT 63.610 2.380 63.780 2.550 ;
        RECT 72.030 3.300 72.200 3.470 ;
        RECT 72.950 3.300 73.120 3.470 ;
        RECT 74.580 3.210 74.750 3.380 ;
        RECT 81.870 3.500 82.040 3.670 ;
        RECT 71.520 2.860 71.690 3.030 ;
        RECT 65.560 2.040 65.730 2.210 ;
        RECT 62.510 1.630 62.680 1.800 ;
        RECT 64.150 1.630 64.320 1.800 ;
        RECT 65.060 1.630 65.230 1.800 ;
        RECT 66.670 1.670 66.840 1.840 ;
        RECT 69.360 2.380 69.530 2.550 ;
        RECT 77.780 3.300 77.950 3.470 ;
        RECT 78.700 3.300 78.870 3.470 ;
        RECT 80.330 3.210 80.500 3.380 ;
        RECT 87.620 3.500 87.790 3.670 ;
        RECT 77.270 2.860 77.440 3.030 ;
        RECT 71.310 2.040 71.480 2.210 ;
        RECT 68.260 1.630 68.430 1.800 ;
        RECT 69.900 1.630 70.070 1.800 ;
        RECT 70.810 1.630 70.980 1.800 ;
        RECT 72.420 1.670 72.590 1.840 ;
        RECT 75.110 2.380 75.280 2.550 ;
        RECT 83.530 3.300 83.700 3.470 ;
        RECT 84.450 3.300 84.620 3.470 ;
        RECT 86.080 3.210 86.250 3.380 ;
        RECT 93.370 3.500 93.540 3.670 ;
        RECT 83.020 2.860 83.190 3.030 ;
        RECT 77.060 2.040 77.230 2.210 ;
        RECT 74.010 1.630 74.180 1.800 ;
        RECT 75.650 1.630 75.820 1.800 ;
        RECT 76.560 1.630 76.730 1.800 ;
        RECT 78.170 1.670 78.340 1.840 ;
        RECT 80.860 2.380 81.030 2.550 ;
        RECT 89.280 3.300 89.450 3.470 ;
        RECT 90.200 3.300 90.370 3.470 ;
        RECT 91.830 3.210 92.000 3.380 ;
        RECT 88.770 2.860 88.940 3.030 ;
        RECT 82.810 2.040 82.980 2.210 ;
        RECT 79.760 1.630 79.930 1.800 ;
        RECT 81.400 1.630 81.570 1.800 ;
        RECT 82.310 1.630 82.480 1.800 ;
        RECT 83.920 1.670 84.090 1.840 ;
        RECT 86.610 2.380 86.780 2.550 ;
        RECT 88.560 2.040 88.730 2.210 ;
        RECT 85.510 1.630 85.680 1.800 ;
        RECT 87.150 1.630 87.320 1.800 ;
        RECT 88.060 1.630 88.230 1.800 ;
        RECT 89.670 1.670 89.840 1.840 ;
        RECT 92.360 2.380 92.530 2.550 ;
        RECT 94.310 2.040 94.480 2.210 ;
        RECT 91.260 1.630 91.430 1.800 ;
        RECT 92.900 1.630 93.070 1.800 ;
        RECT 93.810 1.630 93.980 1.800 ;
        RECT 7.120 1.090 7.290 1.260 ;
        RECT 3.030 0.890 3.200 1.060 ;
        RECT 3.950 0.890 4.120 1.060 ;
        RECT 5.580 0.800 5.750 0.970 ;
        RECT 12.870 1.090 13.040 1.260 ;
        RECT 2.520 0.450 2.690 0.620 ;
        RECT 8.780 0.890 8.950 1.060 ;
        RECT 9.700 0.890 9.870 1.060 ;
        RECT 11.330 0.800 11.500 0.970 ;
        RECT 18.620 1.090 18.790 1.260 ;
        RECT 8.270 0.450 8.440 0.620 ;
        RECT 3.420 -0.740 3.590 -0.570 ;
        RECT 6.110 -0.030 6.280 0.140 ;
        RECT 14.530 0.890 14.700 1.060 ;
        RECT 15.450 0.890 15.620 1.060 ;
        RECT 17.080 0.800 17.250 0.970 ;
        RECT 24.370 1.090 24.540 1.260 ;
        RECT 14.020 0.450 14.190 0.620 ;
        RECT 8.060 -0.370 8.230 -0.200 ;
        RECT 5.010 -0.780 5.180 -0.610 ;
        RECT 6.650 -0.780 6.820 -0.610 ;
        RECT 7.560 -0.780 7.730 -0.610 ;
        RECT 9.170 -0.740 9.340 -0.570 ;
        RECT 11.860 -0.030 12.030 0.140 ;
        RECT 20.280 0.890 20.450 1.060 ;
        RECT 21.200 0.890 21.370 1.060 ;
        RECT 22.830 0.800 23.000 0.970 ;
        RECT 30.120 1.090 30.290 1.260 ;
        RECT 19.770 0.450 19.940 0.620 ;
        RECT 13.810 -0.370 13.980 -0.200 ;
        RECT 10.760 -0.780 10.930 -0.610 ;
        RECT 12.400 -0.780 12.570 -0.610 ;
        RECT 13.310 -0.780 13.480 -0.610 ;
        RECT 14.920 -0.740 15.090 -0.570 ;
        RECT 17.610 -0.030 17.780 0.140 ;
        RECT 26.030 0.890 26.200 1.060 ;
        RECT 26.950 0.890 27.120 1.060 ;
        RECT 28.580 0.800 28.750 0.970 ;
        RECT 35.870 1.090 36.040 1.260 ;
        RECT 25.520 0.450 25.690 0.620 ;
        RECT 19.560 -0.370 19.730 -0.200 ;
        RECT 16.510 -0.780 16.680 -0.610 ;
        RECT 18.150 -0.780 18.320 -0.610 ;
        RECT 19.060 -0.780 19.230 -0.610 ;
        RECT 20.670 -0.740 20.840 -0.570 ;
        RECT 23.360 -0.030 23.530 0.140 ;
        RECT 31.780 0.890 31.950 1.060 ;
        RECT 32.700 0.890 32.870 1.060 ;
        RECT 34.330 0.800 34.500 0.970 ;
        RECT 41.620 1.090 41.790 1.260 ;
        RECT 31.270 0.450 31.440 0.620 ;
        RECT 25.310 -0.370 25.480 -0.200 ;
        RECT 22.260 -0.780 22.430 -0.610 ;
        RECT 23.900 -0.780 24.070 -0.610 ;
        RECT 24.810 -0.780 24.980 -0.610 ;
        RECT 26.420 -0.740 26.590 -0.570 ;
        RECT 29.110 -0.030 29.280 0.140 ;
        RECT 37.530 0.890 37.700 1.060 ;
        RECT 38.450 0.890 38.620 1.060 ;
        RECT 40.080 0.800 40.250 0.970 ;
        RECT 47.370 1.090 47.540 1.260 ;
        RECT 37.020 0.450 37.190 0.620 ;
        RECT 31.060 -0.370 31.230 -0.200 ;
        RECT 28.010 -0.780 28.180 -0.610 ;
        RECT 29.650 -0.780 29.820 -0.610 ;
        RECT 30.560 -0.780 30.730 -0.610 ;
        RECT 32.170 -0.740 32.340 -0.570 ;
        RECT 34.860 -0.030 35.030 0.140 ;
        RECT 43.280 0.890 43.450 1.060 ;
        RECT 44.200 0.890 44.370 1.060 ;
        RECT 45.830 0.800 46.000 0.970 ;
        RECT 53.120 1.090 53.290 1.260 ;
        RECT 42.770 0.450 42.940 0.620 ;
        RECT 36.810 -0.370 36.980 -0.200 ;
        RECT 33.760 -0.780 33.930 -0.610 ;
        RECT 35.400 -0.780 35.570 -0.610 ;
        RECT 36.310 -0.780 36.480 -0.610 ;
        RECT 37.920 -0.740 38.090 -0.570 ;
        RECT 40.610 -0.030 40.780 0.140 ;
        RECT 49.030 0.890 49.200 1.060 ;
        RECT 49.950 0.890 50.120 1.060 ;
        RECT 51.580 0.800 51.750 0.970 ;
        RECT 58.870 1.090 59.040 1.260 ;
        RECT 48.520 0.450 48.690 0.620 ;
        RECT 42.560 -0.370 42.730 -0.200 ;
        RECT 39.510 -0.780 39.680 -0.610 ;
        RECT 41.150 -0.780 41.320 -0.610 ;
        RECT 42.060 -0.780 42.230 -0.610 ;
        RECT 43.670 -0.740 43.840 -0.570 ;
        RECT 46.360 -0.030 46.530 0.140 ;
        RECT 54.780 0.890 54.950 1.060 ;
        RECT 55.700 0.890 55.870 1.060 ;
        RECT 57.330 0.800 57.500 0.970 ;
        RECT 64.620 1.090 64.790 1.260 ;
        RECT 54.270 0.450 54.440 0.620 ;
        RECT 48.310 -0.370 48.480 -0.200 ;
        RECT 45.260 -0.780 45.430 -0.610 ;
        RECT 46.900 -0.780 47.070 -0.610 ;
        RECT 47.810 -0.780 47.980 -0.610 ;
        RECT 49.420 -0.740 49.590 -0.570 ;
        RECT 52.110 -0.030 52.280 0.140 ;
        RECT 60.530 0.890 60.700 1.060 ;
        RECT 61.450 0.890 61.620 1.060 ;
        RECT 63.080 0.800 63.250 0.970 ;
        RECT 70.370 1.090 70.540 1.260 ;
        RECT 60.020 0.450 60.190 0.620 ;
        RECT 54.060 -0.370 54.230 -0.200 ;
        RECT 51.010 -0.780 51.180 -0.610 ;
        RECT 52.650 -0.780 52.820 -0.610 ;
        RECT 53.560 -0.780 53.730 -0.610 ;
        RECT 55.170 -0.740 55.340 -0.570 ;
        RECT 57.860 -0.030 58.030 0.140 ;
        RECT 66.280 0.890 66.450 1.060 ;
        RECT 67.200 0.890 67.370 1.060 ;
        RECT 68.830 0.800 69.000 0.970 ;
        RECT 76.120 1.090 76.290 1.260 ;
        RECT 65.770 0.450 65.940 0.620 ;
        RECT 59.810 -0.370 59.980 -0.200 ;
        RECT 56.760 -0.780 56.930 -0.610 ;
        RECT 58.400 -0.780 58.570 -0.610 ;
        RECT 59.310 -0.780 59.480 -0.610 ;
        RECT 60.920 -0.740 61.090 -0.570 ;
        RECT 63.610 -0.030 63.780 0.140 ;
        RECT 72.030 0.890 72.200 1.060 ;
        RECT 72.950 0.890 73.120 1.060 ;
        RECT 74.580 0.800 74.750 0.970 ;
        RECT 81.870 1.090 82.040 1.260 ;
        RECT 71.520 0.450 71.690 0.620 ;
        RECT 65.560 -0.370 65.730 -0.200 ;
        RECT 62.510 -0.780 62.680 -0.610 ;
        RECT 64.150 -0.780 64.320 -0.610 ;
        RECT 65.060 -0.780 65.230 -0.610 ;
        RECT 66.670 -0.740 66.840 -0.570 ;
        RECT 69.360 -0.030 69.530 0.140 ;
        RECT 77.780 0.890 77.950 1.060 ;
        RECT 78.700 0.890 78.870 1.060 ;
        RECT 80.330 0.800 80.500 0.970 ;
        RECT 87.620 1.090 87.790 1.260 ;
        RECT 77.270 0.450 77.440 0.620 ;
        RECT 71.310 -0.370 71.480 -0.200 ;
        RECT 68.260 -0.780 68.430 -0.610 ;
        RECT 69.900 -0.780 70.070 -0.610 ;
        RECT 70.810 -0.780 70.980 -0.610 ;
        RECT 72.420 -0.740 72.590 -0.570 ;
        RECT 75.110 -0.030 75.280 0.140 ;
        RECT 83.530 0.890 83.700 1.060 ;
        RECT 84.450 0.890 84.620 1.060 ;
        RECT 86.080 0.800 86.250 0.970 ;
        RECT 93.370 1.090 93.540 1.260 ;
        RECT 83.020 0.450 83.190 0.620 ;
        RECT 77.060 -0.370 77.230 -0.200 ;
        RECT 74.010 -0.780 74.180 -0.610 ;
        RECT 75.650 -0.780 75.820 -0.610 ;
        RECT 76.560 -0.780 76.730 -0.610 ;
        RECT 78.170 -0.740 78.340 -0.570 ;
        RECT 80.860 -0.030 81.030 0.140 ;
        RECT 89.280 0.890 89.450 1.060 ;
        RECT 90.200 0.890 90.370 1.060 ;
        RECT 91.830 0.800 92.000 0.970 ;
        RECT 88.770 0.450 88.940 0.620 ;
        RECT 82.810 -0.370 82.980 -0.200 ;
        RECT 79.760 -0.780 79.930 -0.610 ;
        RECT 81.400 -0.780 81.570 -0.610 ;
        RECT 82.310 -0.780 82.480 -0.610 ;
        RECT 83.920 -0.740 84.090 -0.570 ;
        RECT 86.610 -0.030 86.780 0.140 ;
        RECT 88.560 -0.370 88.730 -0.200 ;
        RECT 85.510 -0.780 85.680 -0.610 ;
        RECT 87.150 -0.780 87.320 -0.610 ;
        RECT 88.060 -0.780 88.230 -0.610 ;
        RECT 89.670 -0.740 89.840 -0.570 ;
        RECT 92.360 -0.030 92.530 0.140 ;
        RECT 94.310 -0.370 94.480 -0.200 ;
        RECT 91.260 -0.780 91.430 -0.610 ;
        RECT 92.900 -0.780 93.070 -0.610 ;
        RECT 93.810 -0.780 93.980 -0.610 ;
        RECT 7.120 -1.320 7.290 -1.150 ;
        RECT 3.030 -1.520 3.200 -1.350 ;
        RECT 3.950 -1.520 4.120 -1.350 ;
        RECT 5.580 -1.610 5.750 -1.440 ;
        RECT 12.870 -1.320 13.040 -1.150 ;
        RECT 2.520 -1.960 2.690 -1.790 ;
        RECT 8.780 -1.520 8.950 -1.350 ;
        RECT 9.700 -1.520 9.870 -1.350 ;
        RECT 11.330 -1.610 11.500 -1.440 ;
        RECT 18.620 -1.320 18.790 -1.150 ;
        RECT 8.270 -1.960 8.440 -1.790 ;
        RECT 3.420 -3.150 3.590 -2.980 ;
        RECT 6.110 -2.440 6.280 -2.270 ;
        RECT 14.530 -1.520 14.700 -1.350 ;
        RECT 15.450 -1.520 15.620 -1.350 ;
        RECT 17.080 -1.610 17.250 -1.440 ;
        RECT 24.370 -1.320 24.540 -1.150 ;
        RECT 14.020 -1.960 14.190 -1.790 ;
        RECT 8.060 -2.780 8.230 -2.610 ;
        RECT 5.010 -3.190 5.180 -3.020 ;
        RECT 6.650 -3.190 6.820 -3.020 ;
        RECT 7.560 -3.190 7.730 -3.020 ;
        RECT 9.170 -3.150 9.340 -2.980 ;
        RECT 11.860 -2.440 12.030 -2.270 ;
        RECT 20.280 -1.520 20.450 -1.350 ;
        RECT 21.200 -1.520 21.370 -1.350 ;
        RECT 22.830 -1.610 23.000 -1.440 ;
        RECT 30.120 -1.320 30.290 -1.150 ;
        RECT 19.770 -1.960 19.940 -1.790 ;
        RECT 13.810 -2.780 13.980 -2.610 ;
        RECT 10.760 -3.190 10.930 -3.020 ;
        RECT 12.400 -3.190 12.570 -3.020 ;
        RECT 13.310 -3.190 13.480 -3.020 ;
        RECT 14.920 -3.150 15.090 -2.980 ;
        RECT 17.610 -2.440 17.780 -2.270 ;
        RECT 26.030 -1.520 26.200 -1.350 ;
        RECT 26.950 -1.520 27.120 -1.350 ;
        RECT 28.580 -1.610 28.750 -1.440 ;
        RECT 35.870 -1.320 36.040 -1.150 ;
        RECT 25.520 -1.960 25.690 -1.790 ;
        RECT 19.560 -2.780 19.730 -2.610 ;
        RECT 16.510 -3.190 16.680 -3.020 ;
        RECT 18.150 -3.190 18.320 -3.020 ;
        RECT 19.060 -3.190 19.230 -3.020 ;
        RECT 20.670 -3.150 20.840 -2.980 ;
        RECT 23.360 -2.440 23.530 -2.270 ;
        RECT 31.780 -1.520 31.950 -1.350 ;
        RECT 32.700 -1.520 32.870 -1.350 ;
        RECT 34.330 -1.610 34.500 -1.440 ;
        RECT 41.620 -1.320 41.790 -1.150 ;
        RECT 31.270 -1.960 31.440 -1.790 ;
        RECT 25.310 -2.780 25.480 -2.610 ;
        RECT 22.260 -3.190 22.430 -3.020 ;
        RECT 23.900 -3.190 24.070 -3.020 ;
        RECT 24.810 -3.190 24.980 -3.020 ;
        RECT 26.420 -3.150 26.590 -2.980 ;
        RECT 29.110 -2.440 29.280 -2.270 ;
        RECT 37.530 -1.520 37.700 -1.350 ;
        RECT 38.450 -1.520 38.620 -1.350 ;
        RECT 40.080 -1.610 40.250 -1.440 ;
        RECT 47.370 -1.320 47.540 -1.150 ;
        RECT 37.020 -1.960 37.190 -1.790 ;
        RECT 31.060 -2.780 31.230 -2.610 ;
        RECT 28.010 -3.190 28.180 -3.020 ;
        RECT 29.650 -3.190 29.820 -3.020 ;
        RECT 30.560 -3.190 30.730 -3.020 ;
        RECT 32.170 -3.150 32.340 -2.980 ;
        RECT 34.860 -2.440 35.030 -2.270 ;
        RECT 43.280 -1.520 43.450 -1.350 ;
        RECT 44.200 -1.520 44.370 -1.350 ;
        RECT 45.830 -1.610 46.000 -1.440 ;
        RECT 53.120 -1.320 53.290 -1.150 ;
        RECT 42.770 -1.960 42.940 -1.790 ;
        RECT 36.810 -2.780 36.980 -2.610 ;
        RECT 33.760 -3.190 33.930 -3.020 ;
        RECT 35.400 -3.190 35.570 -3.020 ;
        RECT 36.310 -3.190 36.480 -3.020 ;
        RECT 37.920 -3.150 38.090 -2.980 ;
        RECT 40.610 -2.440 40.780 -2.270 ;
        RECT 49.030 -1.520 49.200 -1.350 ;
        RECT 49.950 -1.520 50.120 -1.350 ;
        RECT 51.580 -1.610 51.750 -1.440 ;
        RECT 58.870 -1.320 59.040 -1.150 ;
        RECT 48.520 -1.960 48.690 -1.790 ;
        RECT 42.560 -2.780 42.730 -2.610 ;
        RECT 39.510 -3.190 39.680 -3.020 ;
        RECT 41.150 -3.190 41.320 -3.020 ;
        RECT 42.060 -3.190 42.230 -3.020 ;
        RECT 43.670 -3.150 43.840 -2.980 ;
        RECT 46.360 -2.440 46.530 -2.270 ;
        RECT 54.780 -1.520 54.950 -1.350 ;
        RECT 55.700 -1.520 55.870 -1.350 ;
        RECT 57.330 -1.610 57.500 -1.440 ;
        RECT 64.620 -1.320 64.790 -1.150 ;
        RECT 54.270 -1.960 54.440 -1.790 ;
        RECT 48.310 -2.780 48.480 -2.610 ;
        RECT 45.260 -3.190 45.430 -3.020 ;
        RECT 46.900 -3.190 47.070 -3.020 ;
        RECT 47.810 -3.190 47.980 -3.020 ;
        RECT 49.420 -3.150 49.590 -2.980 ;
        RECT 52.110 -2.440 52.280 -2.270 ;
        RECT 60.530 -1.520 60.700 -1.350 ;
        RECT 61.450 -1.520 61.620 -1.350 ;
        RECT 63.080 -1.610 63.250 -1.440 ;
        RECT 70.370 -1.320 70.540 -1.150 ;
        RECT 60.020 -1.960 60.190 -1.790 ;
        RECT 54.060 -2.780 54.230 -2.610 ;
        RECT 51.010 -3.190 51.180 -3.020 ;
        RECT 52.650 -3.190 52.820 -3.020 ;
        RECT 53.560 -3.190 53.730 -3.020 ;
        RECT 55.170 -3.150 55.340 -2.980 ;
        RECT 57.860 -2.440 58.030 -2.270 ;
        RECT 66.280 -1.520 66.450 -1.350 ;
        RECT 67.200 -1.520 67.370 -1.350 ;
        RECT 68.830 -1.610 69.000 -1.440 ;
        RECT 76.120 -1.320 76.290 -1.150 ;
        RECT 65.770 -1.960 65.940 -1.790 ;
        RECT 59.810 -2.780 59.980 -2.610 ;
        RECT 56.760 -3.190 56.930 -3.020 ;
        RECT 58.400 -3.190 58.570 -3.020 ;
        RECT 59.310 -3.190 59.480 -3.020 ;
        RECT 60.920 -3.150 61.090 -2.980 ;
        RECT 63.610 -2.440 63.780 -2.270 ;
        RECT 72.030 -1.520 72.200 -1.350 ;
        RECT 72.950 -1.520 73.120 -1.350 ;
        RECT 74.580 -1.610 74.750 -1.440 ;
        RECT 81.870 -1.320 82.040 -1.150 ;
        RECT 71.520 -1.960 71.690 -1.790 ;
        RECT 65.560 -2.780 65.730 -2.610 ;
        RECT 62.510 -3.190 62.680 -3.020 ;
        RECT 64.150 -3.190 64.320 -3.020 ;
        RECT 65.060 -3.190 65.230 -3.020 ;
        RECT 66.670 -3.150 66.840 -2.980 ;
        RECT 69.360 -2.440 69.530 -2.270 ;
        RECT 77.780 -1.520 77.950 -1.350 ;
        RECT 78.700 -1.520 78.870 -1.350 ;
        RECT 80.330 -1.610 80.500 -1.440 ;
        RECT 87.620 -1.320 87.790 -1.150 ;
        RECT 77.270 -1.960 77.440 -1.790 ;
        RECT 71.310 -2.780 71.480 -2.610 ;
        RECT 68.260 -3.190 68.430 -3.020 ;
        RECT 69.900 -3.190 70.070 -3.020 ;
        RECT 70.810 -3.190 70.980 -3.020 ;
        RECT 72.420 -3.150 72.590 -2.980 ;
        RECT 75.110 -2.440 75.280 -2.270 ;
        RECT 83.530 -1.520 83.700 -1.350 ;
        RECT 84.450 -1.520 84.620 -1.350 ;
        RECT 86.080 -1.610 86.250 -1.440 ;
        RECT 93.370 -1.320 93.540 -1.150 ;
        RECT 83.020 -1.960 83.190 -1.790 ;
        RECT 77.060 -2.780 77.230 -2.610 ;
        RECT 74.010 -3.190 74.180 -3.020 ;
        RECT 75.650 -3.190 75.820 -3.020 ;
        RECT 76.560 -3.190 76.730 -3.020 ;
        RECT 78.170 -3.150 78.340 -2.980 ;
        RECT 80.860 -2.440 81.030 -2.270 ;
        RECT 89.280 -1.520 89.450 -1.350 ;
        RECT 90.200 -1.520 90.370 -1.350 ;
        RECT 91.830 -1.610 92.000 -1.440 ;
        RECT 88.770 -1.960 88.940 -1.790 ;
        RECT 82.810 -2.780 82.980 -2.610 ;
        RECT 79.760 -3.190 79.930 -3.020 ;
        RECT 81.400 -3.190 81.570 -3.020 ;
        RECT 82.310 -3.190 82.480 -3.020 ;
        RECT 83.920 -3.150 84.090 -2.980 ;
        RECT 86.610 -2.440 86.780 -2.270 ;
        RECT 88.560 -2.780 88.730 -2.610 ;
        RECT 85.510 -3.190 85.680 -3.020 ;
        RECT 87.150 -3.190 87.320 -3.020 ;
        RECT 88.060 -3.190 88.230 -3.020 ;
        RECT 89.670 -3.150 89.840 -2.980 ;
        RECT 92.360 -2.440 92.530 -2.270 ;
        RECT 94.310 -2.780 94.480 -2.610 ;
        RECT 91.260 -3.190 91.430 -3.020 ;
        RECT 92.900 -3.190 93.070 -3.020 ;
        RECT 93.810 -3.190 93.980 -3.020 ;
        RECT 7.120 -3.730 7.290 -3.560 ;
        RECT 3.030 -3.930 3.200 -3.760 ;
        RECT 3.950 -3.930 4.120 -3.760 ;
        RECT 5.580 -4.020 5.750 -3.850 ;
        RECT 12.870 -3.730 13.040 -3.560 ;
        RECT 2.520 -4.370 2.690 -4.200 ;
        RECT 8.780 -3.930 8.950 -3.760 ;
        RECT 9.700 -3.930 9.870 -3.760 ;
        RECT 11.330 -4.020 11.500 -3.850 ;
        RECT 18.620 -3.730 18.790 -3.560 ;
        RECT 8.270 -4.370 8.440 -4.200 ;
        RECT 3.420 -5.560 3.590 -5.390 ;
        RECT 6.110 -4.850 6.280 -4.680 ;
        RECT 14.530 -3.930 14.700 -3.760 ;
        RECT 15.450 -3.930 15.620 -3.760 ;
        RECT 17.080 -4.020 17.250 -3.850 ;
        RECT 24.370 -3.730 24.540 -3.560 ;
        RECT 14.020 -4.370 14.190 -4.200 ;
        RECT 8.060 -5.190 8.230 -5.020 ;
        RECT 5.010 -5.600 5.180 -5.430 ;
        RECT 6.650 -5.600 6.820 -5.430 ;
        RECT 7.560 -5.600 7.730 -5.430 ;
        RECT 7.120 -6.460 7.290 -6.290 ;
        RECT 9.170 -5.560 9.340 -5.390 ;
        RECT 11.860 -4.850 12.030 -4.680 ;
        RECT 20.280 -3.930 20.450 -3.760 ;
        RECT 21.200 -3.930 21.370 -3.760 ;
        RECT 22.830 -4.020 23.000 -3.850 ;
        RECT 30.120 -3.730 30.290 -3.560 ;
        RECT 19.770 -4.370 19.940 -4.200 ;
        RECT 13.810 -5.190 13.980 -5.020 ;
        RECT 10.760 -5.600 10.930 -5.430 ;
        RECT 12.400 -5.600 12.570 -5.430 ;
        RECT 13.310 -5.600 13.480 -5.430 ;
        RECT 3.030 -6.930 3.200 -6.760 ;
        RECT 3.950 -6.930 4.120 -6.760 ;
        RECT 5.580 -7.020 5.750 -6.850 ;
        RECT 12.870 -6.460 13.040 -6.290 ;
        RECT 14.920 -5.560 15.090 -5.390 ;
        RECT 17.610 -4.850 17.780 -4.680 ;
        RECT 26.030 -3.930 26.200 -3.760 ;
        RECT 26.950 -3.930 27.120 -3.760 ;
        RECT 28.580 -4.020 28.750 -3.850 ;
        RECT 35.870 -3.730 36.040 -3.560 ;
        RECT 25.520 -4.370 25.690 -4.200 ;
        RECT 19.560 -5.190 19.730 -5.020 ;
        RECT 16.510 -5.600 16.680 -5.430 ;
        RECT 18.150 -5.600 18.320 -5.430 ;
        RECT 19.060 -5.600 19.230 -5.430 ;
        RECT 2.520 -7.370 2.690 -7.200 ;
        RECT 8.780 -6.930 8.950 -6.760 ;
        RECT 9.700 -6.930 9.870 -6.760 ;
        RECT 11.330 -7.020 11.500 -6.850 ;
        RECT 18.620 -6.460 18.790 -6.290 ;
        RECT 20.670 -5.560 20.840 -5.390 ;
        RECT 23.360 -4.850 23.530 -4.680 ;
        RECT 31.780 -3.930 31.950 -3.760 ;
        RECT 32.700 -3.930 32.870 -3.760 ;
        RECT 34.330 -4.020 34.500 -3.850 ;
        RECT 41.620 -3.730 41.790 -3.560 ;
        RECT 31.270 -4.370 31.440 -4.200 ;
        RECT 25.310 -5.190 25.480 -5.020 ;
        RECT 22.260 -5.600 22.430 -5.430 ;
        RECT 23.900 -5.600 24.070 -5.430 ;
        RECT 24.810 -5.600 24.980 -5.430 ;
        RECT 8.270 -7.370 8.440 -7.200 ;
        RECT 3.420 -8.560 3.590 -8.390 ;
        RECT 6.110 -7.850 6.280 -7.680 ;
        RECT 14.530 -6.930 14.700 -6.760 ;
        RECT 15.450 -6.930 15.620 -6.760 ;
        RECT 17.080 -7.020 17.250 -6.850 ;
        RECT 24.370 -6.460 24.540 -6.290 ;
        RECT 26.420 -5.560 26.590 -5.390 ;
        RECT 29.110 -4.850 29.280 -4.680 ;
        RECT 37.530 -3.930 37.700 -3.760 ;
        RECT 38.450 -3.930 38.620 -3.760 ;
        RECT 40.080 -4.020 40.250 -3.850 ;
        RECT 47.370 -3.730 47.540 -3.560 ;
        RECT 37.020 -4.370 37.190 -4.200 ;
        RECT 31.060 -5.190 31.230 -5.020 ;
        RECT 28.010 -5.600 28.180 -5.430 ;
        RECT 29.650 -5.600 29.820 -5.430 ;
        RECT 30.560 -5.600 30.730 -5.430 ;
        RECT 14.020 -7.370 14.190 -7.200 ;
        RECT 8.060 -8.190 8.230 -8.020 ;
        RECT 5.010 -8.600 5.180 -8.430 ;
        RECT 6.650 -8.600 6.820 -8.430 ;
        RECT 7.560 -8.600 7.730 -8.430 ;
        RECT 9.170 -8.560 9.340 -8.390 ;
        RECT 11.860 -7.850 12.030 -7.680 ;
        RECT 20.280 -6.930 20.450 -6.760 ;
        RECT 21.200 -6.930 21.370 -6.760 ;
        RECT 22.830 -7.020 23.000 -6.850 ;
        RECT 30.120 -6.460 30.290 -6.290 ;
        RECT 32.170 -5.560 32.340 -5.390 ;
        RECT 34.860 -4.850 35.030 -4.680 ;
        RECT 43.280 -3.930 43.450 -3.760 ;
        RECT 44.200 -3.930 44.370 -3.760 ;
        RECT 45.830 -4.020 46.000 -3.850 ;
        RECT 53.120 -3.730 53.290 -3.560 ;
        RECT 42.770 -4.370 42.940 -4.200 ;
        RECT 36.810 -5.190 36.980 -5.020 ;
        RECT 33.760 -5.600 33.930 -5.430 ;
        RECT 35.400 -5.600 35.570 -5.430 ;
        RECT 36.310 -5.600 36.480 -5.430 ;
        RECT 19.770 -7.370 19.940 -7.200 ;
        RECT 13.810 -8.190 13.980 -8.020 ;
        RECT 10.760 -8.600 10.930 -8.430 ;
        RECT 12.400 -8.600 12.570 -8.430 ;
        RECT 13.310 -8.600 13.480 -8.430 ;
        RECT 14.920 -8.560 15.090 -8.390 ;
        RECT 17.610 -7.850 17.780 -7.680 ;
        RECT 26.030 -6.930 26.200 -6.760 ;
        RECT 26.950 -6.930 27.120 -6.760 ;
        RECT 28.580 -7.020 28.750 -6.850 ;
        RECT 35.870 -6.460 36.040 -6.290 ;
        RECT 37.920 -5.560 38.090 -5.390 ;
        RECT 40.610 -4.850 40.780 -4.680 ;
        RECT 49.030 -3.930 49.200 -3.760 ;
        RECT 49.950 -3.930 50.120 -3.760 ;
        RECT 51.580 -4.020 51.750 -3.850 ;
        RECT 58.870 -3.730 59.040 -3.560 ;
        RECT 48.520 -4.370 48.690 -4.200 ;
        RECT 42.560 -5.190 42.730 -5.020 ;
        RECT 39.510 -5.600 39.680 -5.430 ;
        RECT 41.150 -5.600 41.320 -5.430 ;
        RECT 42.060 -5.600 42.230 -5.430 ;
        RECT 25.520 -7.370 25.690 -7.200 ;
        RECT 19.560 -8.190 19.730 -8.020 ;
        RECT 16.510 -8.600 16.680 -8.430 ;
        RECT 18.150 -8.600 18.320 -8.430 ;
        RECT 19.060 -8.600 19.230 -8.430 ;
        RECT 20.670 -8.560 20.840 -8.390 ;
        RECT 23.360 -7.850 23.530 -7.680 ;
        RECT 31.780 -6.930 31.950 -6.760 ;
        RECT 32.700 -6.930 32.870 -6.760 ;
        RECT 34.330 -7.020 34.500 -6.850 ;
        RECT 41.620 -6.460 41.790 -6.290 ;
        RECT 43.670 -5.560 43.840 -5.390 ;
        RECT 46.360 -4.850 46.530 -4.680 ;
        RECT 54.780 -3.930 54.950 -3.760 ;
        RECT 55.700 -3.930 55.870 -3.760 ;
        RECT 57.330 -4.020 57.500 -3.850 ;
        RECT 64.620 -3.730 64.790 -3.560 ;
        RECT 54.270 -4.370 54.440 -4.200 ;
        RECT 48.310 -5.190 48.480 -5.020 ;
        RECT 45.260 -5.600 45.430 -5.430 ;
        RECT 46.900 -5.600 47.070 -5.430 ;
        RECT 47.810 -5.600 47.980 -5.430 ;
        RECT 31.270 -7.370 31.440 -7.200 ;
        RECT 25.310 -8.190 25.480 -8.020 ;
        RECT 22.260 -8.600 22.430 -8.430 ;
        RECT 23.900 -8.600 24.070 -8.430 ;
        RECT 24.810 -8.600 24.980 -8.430 ;
        RECT 26.420 -8.560 26.590 -8.390 ;
        RECT 29.110 -7.850 29.280 -7.680 ;
        RECT 37.530 -6.930 37.700 -6.760 ;
        RECT 38.450 -6.930 38.620 -6.760 ;
        RECT 40.080 -7.020 40.250 -6.850 ;
        RECT 47.370 -6.460 47.540 -6.290 ;
        RECT 49.420 -5.560 49.590 -5.390 ;
        RECT 52.110 -4.850 52.280 -4.680 ;
        RECT 60.530 -3.930 60.700 -3.760 ;
        RECT 61.450 -3.930 61.620 -3.760 ;
        RECT 63.080 -4.020 63.250 -3.850 ;
        RECT 70.370 -3.730 70.540 -3.560 ;
        RECT 60.020 -4.370 60.190 -4.200 ;
        RECT 54.060 -5.190 54.230 -5.020 ;
        RECT 51.010 -5.600 51.180 -5.430 ;
        RECT 52.650 -5.600 52.820 -5.430 ;
        RECT 53.560 -5.600 53.730 -5.430 ;
        RECT 37.020 -7.370 37.190 -7.200 ;
        RECT 31.060 -8.190 31.230 -8.020 ;
        RECT 28.010 -8.600 28.180 -8.430 ;
        RECT 29.650 -8.600 29.820 -8.430 ;
        RECT 30.560 -8.600 30.730 -8.430 ;
        RECT 32.170 -8.560 32.340 -8.390 ;
        RECT 34.860 -7.850 35.030 -7.680 ;
        RECT 43.280 -6.930 43.450 -6.760 ;
        RECT 44.200 -6.930 44.370 -6.760 ;
        RECT 45.830 -7.020 46.000 -6.850 ;
        RECT 53.120 -6.460 53.290 -6.290 ;
        RECT 55.170 -5.560 55.340 -5.390 ;
        RECT 57.860 -4.850 58.030 -4.680 ;
        RECT 66.280 -3.930 66.450 -3.760 ;
        RECT 67.200 -3.930 67.370 -3.760 ;
        RECT 68.830 -4.020 69.000 -3.850 ;
        RECT 76.120 -3.730 76.290 -3.560 ;
        RECT 65.770 -4.370 65.940 -4.200 ;
        RECT 59.810 -5.190 59.980 -5.020 ;
        RECT 56.760 -5.600 56.930 -5.430 ;
        RECT 58.400 -5.600 58.570 -5.430 ;
        RECT 59.310 -5.600 59.480 -5.430 ;
        RECT 42.770 -7.370 42.940 -7.200 ;
        RECT 36.810 -8.190 36.980 -8.020 ;
        RECT 33.760 -8.600 33.930 -8.430 ;
        RECT 35.400 -8.600 35.570 -8.430 ;
        RECT 36.310 -8.600 36.480 -8.430 ;
        RECT 37.920 -8.560 38.090 -8.390 ;
        RECT 40.610 -7.850 40.780 -7.680 ;
        RECT 49.030 -6.930 49.200 -6.760 ;
        RECT 49.950 -6.930 50.120 -6.760 ;
        RECT 51.580 -7.020 51.750 -6.850 ;
        RECT 58.870 -6.460 59.040 -6.290 ;
        RECT 60.920 -5.560 61.090 -5.390 ;
        RECT 63.610 -4.850 63.780 -4.680 ;
        RECT 72.030 -3.930 72.200 -3.760 ;
        RECT 72.950 -3.930 73.120 -3.760 ;
        RECT 74.580 -4.020 74.750 -3.850 ;
        RECT 81.870 -3.730 82.040 -3.560 ;
        RECT 71.520 -4.370 71.690 -4.200 ;
        RECT 65.560 -5.190 65.730 -5.020 ;
        RECT 62.510 -5.600 62.680 -5.430 ;
        RECT 64.150 -5.600 64.320 -5.430 ;
        RECT 65.060 -5.600 65.230 -5.430 ;
        RECT 48.520 -7.370 48.690 -7.200 ;
        RECT 42.560 -8.190 42.730 -8.020 ;
        RECT 39.510 -8.600 39.680 -8.430 ;
        RECT 41.150 -8.600 41.320 -8.430 ;
        RECT 42.060 -8.600 42.230 -8.430 ;
        RECT 43.670 -8.560 43.840 -8.390 ;
        RECT 46.360 -7.850 46.530 -7.680 ;
        RECT 54.780 -6.930 54.950 -6.760 ;
        RECT 55.700 -6.930 55.870 -6.760 ;
        RECT 57.330 -7.020 57.500 -6.850 ;
        RECT 64.620 -6.460 64.790 -6.290 ;
        RECT 66.670 -5.560 66.840 -5.390 ;
        RECT 69.360 -4.850 69.530 -4.680 ;
        RECT 77.780 -3.930 77.950 -3.760 ;
        RECT 78.700 -3.930 78.870 -3.760 ;
        RECT 80.330 -4.020 80.500 -3.850 ;
        RECT 87.620 -3.730 87.790 -3.560 ;
        RECT 77.270 -4.370 77.440 -4.200 ;
        RECT 71.310 -5.190 71.480 -5.020 ;
        RECT 68.260 -5.600 68.430 -5.430 ;
        RECT 69.900 -5.600 70.070 -5.430 ;
        RECT 70.810 -5.600 70.980 -5.430 ;
        RECT 54.270 -7.370 54.440 -7.200 ;
        RECT 48.310 -8.190 48.480 -8.020 ;
        RECT 45.260 -8.600 45.430 -8.430 ;
        RECT 46.900 -8.600 47.070 -8.430 ;
        RECT 47.810 -8.600 47.980 -8.430 ;
        RECT 49.420 -8.560 49.590 -8.390 ;
        RECT 52.110 -7.850 52.280 -7.680 ;
        RECT 60.530 -6.930 60.700 -6.760 ;
        RECT 61.450 -6.930 61.620 -6.760 ;
        RECT 63.080 -7.020 63.250 -6.850 ;
        RECT 70.370 -6.460 70.540 -6.290 ;
        RECT 72.420 -5.560 72.590 -5.390 ;
        RECT 75.110 -4.850 75.280 -4.680 ;
        RECT 83.530 -3.930 83.700 -3.760 ;
        RECT 84.450 -3.930 84.620 -3.760 ;
        RECT 86.080 -4.020 86.250 -3.850 ;
        RECT 93.370 -3.730 93.540 -3.560 ;
        RECT 83.020 -4.370 83.190 -4.200 ;
        RECT 77.060 -5.190 77.230 -5.020 ;
        RECT 74.010 -5.600 74.180 -5.430 ;
        RECT 75.650 -5.600 75.820 -5.430 ;
        RECT 76.560 -5.600 76.730 -5.430 ;
        RECT 60.020 -7.370 60.190 -7.200 ;
        RECT 54.060 -8.190 54.230 -8.020 ;
        RECT 51.010 -8.600 51.180 -8.430 ;
        RECT 52.650 -8.600 52.820 -8.430 ;
        RECT 53.560 -8.600 53.730 -8.430 ;
        RECT 55.170 -8.560 55.340 -8.390 ;
        RECT 57.860 -7.850 58.030 -7.680 ;
        RECT 66.280 -6.930 66.450 -6.760 ;
        RECT 67.200 -6.930 67.370 -6.760 ;
        RECT 68.830 -7.020 69.000 -6.850 ;
        RECT 76.120 -6.460 76.290 -6.290 ;
        RECT 78.170 -5.560 78.340 -5.390 ;
        RECT 80.860 -4.850 81.030 -4.680 ;
        RECT 89.280 -3.930 89.450 -3.760 ;
        RECT 90.200 -3.930 90.370 -3.760 ;
        RECT 91.830 -4.020 92.000 -3.850 ;
        RECT 88.770 -4.370 88.940 -4.200 ;
        RECT 82.810 -5.190 82.980 -5.020 ;
        RECT 79.760 -5.600 79.930 -5.430 ;
        RECT 81.400 -5.600 81.570 -5.430 ;
        RECT 82.310 -5.600 82.480 -5.430 ;
        RECT 65.770 -7.370 65.940 -7.200 ;
        RECT 59.810 -8.190 59.980 -8.020 ;
        RECT 56.760 -8.600 56.930 -8.430 ;
        RECT 58.400 -8.600 58.570 -8.430 ;
        RECT 59.310 -8.600 59.480 -8.430 ;
        RECT 60.920 -8.560 61.090 -8.390 ;
        RECT 63.610 -7.850 63.780 -7.680 ;
        RECT 72.030 -6.930 72.200 -6.760 ;
        RECT 72.950 -6.930 73.120 -6.760 ;
        RECT 74.580 -7.020 74.750 -6.850 ;
        RECT 81.870 -6.460 82.040 -6.290 ;
        RECT 83.920 -5.560 84.090 -5.390 ;
        RECT 86.610 -4.850 86.780 -4.680 ;
        RECT 88.560 -5.190 88.730 -5.020 ;
        RECT 85.510 -5.600 85.680 -5.430 ;
        RECT 87.150 -5.600 87.320 -5.430 ;
        RECT 88.060 -5.600 88.230 -5.430 ;
        RECT 71.520 -7.370 71.690 -7.200 ;
        RECT 65.560 -8.190 65.730 -8.020 ;
        RECT 62.510 -8.600 62.680 -8.430 ;
        RECT 64.150 -8.600 64.320 -8.430 ;
        RECT 65.060 -8.600 65.230 -8.430 ;
        RECT 66.670 -8.560 66.840 -8.390 ;
        RECT 69.360 -7.850 69.530 -7.680 ;
        RECT 77.780 -6.930 77.950 -6.760 ;
        RECT 78.700 -6.930 78.870 -6.760 ;
        RECT 80.330 -7.020 80.500 -6.850 ;
        RECT 87.620 -6.460 87.790 -6.290 ;
        RECT 89.670 -5.560 89.840 -5.390 ;
        RECT 92.360 -4.850 92.530 -4.680 ;
        RECT 94.310 -5.190 94.480 -5.020 ;
        RECT 91.260 -5.600 91.430 -5.430 ;
        RECT 92.900 -5.600 93.070 -5.430 ;
        RECT 93.810 -5.600 93.980 -5.430 ;
        RECT 77.270 -7.370 77.440 -7.200 ;
        RECT 71.310 -8.190 71.480 -8.020 ;
        RECT 68.260 -8.600 68.430 -8.430 ;
        RECT 69.900 -8.600 70.070 -8.430 ;
        RECT 70.810 -8.600 70.980 -8.430 ;
        RECT 72.420 -8.560 72.590 -8.390 ;
        RECT 75.110 -7.850 75.280 -7.680 ;
        RECT 83.530 -6.930 83.700 -6.760 ;
        RECT 84.450 -6.930 84.620 -6.760 ;
        RECT 86.080 -7.020 86.250 -6.850 ;
        RECT 83.020 -7.370 83.190 -7.200 ;
        RECT 77.060 -8.190 77.230 -8.020 ;
        RECT 74.010 -8.600 74.180 -8.430 ;
        RECT 75.650 -8.600 75.820 -8.430 ;
        RECT 76.560 -8.600 76.730 -8.430 ;
        RECT 78.170 -8.560 78.340 -8.390 ;
        RECT 80.860 -7.850 81.030 -7.680 ;
        RECT 89.280 -6.930 89.450 -6.760 ;
        RECT 90.200 -6.930 90.370 -6.760 ;
        RECT 91.830 -7.020 92.000 -6.850 ;
        RECT 88.770 -7.370 88.940 -7.200 ;
        RECT 82.810 -8.190 82.980 -8.020 ;
        RECT 79.760 -8.600 79.930 -8.430 ;
        RECT 81.400 -8.600 81.570 -8.430 ;
        RECT 82.310 -8.600 82.480 -8.430 ;
        RECT 83.920 -8.560 84.090 -8.390 ;
        RECT 86.610 -7.850 86.780 -7.680 ;
        RECT 88.560 -8.190 88.730 -8.020 ;
        RECT 85.510 -8.600 85.680 -8.430 ;
        RECT 87.150 -8.600 87.320 -8.430 ;
        RECT 88.060 -8.600 88.230 -8.430 ;
        RECT 89.670 -8.560 89.840 -8.390 ;
        RECT 92.360 -7.850 92.530 -7.680 ;
        RECT 94.310 -8.190 94.480 -8.020 ;
        RECT 91.260 -8.600 91.430 -8.430 ;
        RECT 92.900 -8.600 93.070 -8.430 ;
        RECT 93.810 -8.600 93.980 -8.430 ;
        RECT 7.120 -9.140 7.290 -8.970 ;
        RECT 3.030 -9.340 3.200 -9.170 ;
        RECT 3.950 -9.340 4.120 -9.170 ;
        RECT 5.580 -9.430 5.750 -9.260 ;
        RECT 12.870 -9.140 13.040 -8.970 ;
        RECT 2.520 -9.780 2.690 -9.610 ;
        RECT 8.780 -9.340 8.950 -9.170 ;
        RECT 9.700 -9.340 9.870 -9.170 ;
        RECT 11.330 -9.430 11.500 -9.260 ;
        RECT 18.620 -9.140 18.790 -8.970 ;
        RECT 8.270 -9.780 8.440 -9.610 ;
        RECT 3.420 -10.970 3.590 -10.800 ;
        RECT 6.110 -10.260 6.280 -10.090 ;
        RECT 14.530 -9.340 14.700 -9.170 ;
        RECT 15.450 -9.340 15.620 -9.170 ;
        RECT 17.080 -9.430 17.250 -9.260 ;
        RECT 24.370 -9.140 24.540 -8.970 ;
        RECT 14.020 -9.780 14.190 -9.610 ;
        RECT 8.060 -10.600 8.230 -10.430 ;
        RECT 5.010 -11.010 5.180 -10.840 ;
        RECT 6.650 -11.010 6.820 -10.840 ;
        RECT 7.560 -11.010 7.730 -10.840 ;
        RECT 9.170 -10.970 9.340 -10.800 ;
        RECT 11.860 -10.260 12.030 -10.090 ;
        RECT 20.280 -9.340 20.450 -9.170 ;
        RECT 21.200 -9.340 21.370 -9.170 ;
        RECT 22.830 -9.430 23.000 -9.260 ;
        RECT 30.120 -9.140 30.290 -8.970 ;
        RECT 19.770 -9.780 19.940 -9.610 ;
        RECT 13.810 -10.600 13.980 -10.430 ;
        RECT 10.760 -11.010 10.930 -10.840 ;
        RECT 12.400 -11.010 12.570 -10.840 ;
        RECT 13.310 -11.010 13.480 -10.840 ;
        RECT 14.920 -10.970 15.090 -10.800 ;
        RECT 17.610 -10.260 17.780 -10.090 ;
        RECT 26.030 -9.340 26.200 -9.170 ;
        RECT 26.950 -9.340 27.120 -9.170 ;
        RECT 28.580 -9.430 28.750 -9.260 ;
        RECT 35.870 -9.140 36.040 -8.970 ;
        RECT 25.520 -9.780 25.690 -9.610 ;
        RECT 19.560 -10.600 19.730 -10.430 ;
        RECT 16.510 -11.010 16.680 -10.840 ;
        RECT 18.150 -11.010 18.320 -10.840 ;
        RECT 19.060 -11.010 19.230 -10.840 ;
        RECT 20.670 -10.970 20.840 -10.800 ;
        RECT 23.360 -10.260 23.530 -10.090 ;
        RECT 31.780 -9.340 31.950 -9.170 ;
        RECT 32.700 -9.340 32.870 -9.170 ;
        RECT 34.330 -9.430 34.500 -9.260 ;
        RECT 41.620 -9.140 41.790 -8.970 ;
        RECT 31.270 -9.780 31.440 -9.610 ;
        RECT 25.310 -10.600 25.480 -10.430 ;
        RECT 22.260 -11.010 22.430 -10.840 ;
        RECT 23.900 -11.010 24.070 -10.840 ;
        RECT 24.810 -11.010 24.980 -10.840 ;
        RECT 26.420 -10.970 26.590 -10.800 ;
        RECT 29.110 -10.260 29.280 -10.090 ;
        RECT 37.530 -9.340 37.700 -9.170 ;
        RECT 38.450 -9.340 38.620 -9.170 ;
        RECT 40.080 -9.430 40.250 -9.260 ;
        RECT 47.370 -9.140 47.540 -8.970 ;
        RECT 37.020 -9.780 37.190 -9.610 ;
        RECT 31.060 -10.600 31.230 -10.430 ;
        RECT 28.010 -11.010 28.180 -10.840 ;
        RECT 29.650 -11.010 29.820 -10.840 ;
        RECT 30.560 -11.010 30.730 -10.840 ;
        RECT 32.170 -10.970 32.340 -10.800 ;
        RECT 34.860 -10.260 35.030 -10.090 ;
        RECT 43.280 -9.340 43.450 -9.170 ;
        RECT 44.200 -9.340 44.370 -9.170 ;
        RECT 45.830 -9.430 46.000 -9.260 ;
        RECT 53.120 -9.140 53.290 -8.970 ;
        RECT 42.770 -9.780 42.940 -9.610 ;
        RECT 36.810 -10.600 36.980 -10.430 ;
        RECT 33.760 -11.010 33.930 -10.840 ;
        RECT 35.400 -11.010 35.570 -10.840 ;
        RECT 36.310 -11.010 36.480 -10.840 ;
        RECT 37.920 -10.970 38.090 -10.800 ;
        RECT 40.610 -10.260 40.780 -10.090 ;
        RECT 49.030 -9.340 49.200 -9.170 ;
        RECT 49.950 -9.340 50.120 -9.170 ;
        RECT 51.580 -9.430 51.750 -9.260 ;
        RECT 58.870 -9.140 59.040 -8.970 ;
        RECT 48.520 -9.780 48.690 -9.610 ;
        RECT 42.560 -10.600 42.730 -10.430 ;
        RECT 39.510 -11.010 39.680 -10.840 ;
        RECT 41.150 -11.010 41.320 -10.840 ;
        RECT 42.060 -11.010 42.230 -10.840 ;
        RECT 43.670 -10.970 43.840 -10.800 ;
        RECT 46.360 -10.260 46.530 -10.090 ;
        RECT 54.780 -9.340 54.950 -9.170 ;
        RECT 55.700 -9.340 55.870 -9.170 ;
        RECT 57.330 -9.430 57.500 -9.260 ;
        RECT 64.620 -9.140 64.790 -8.970 ;
        RECT 54.270 -9.780 54.440 -9.610 ;
        RECT 48.310 -10.600 48.480 -10.430 ;
        RECT 45.260 -11.010 45.430 -10.840 ;
        RECT 46.900 -11.010 47.070 -10.840 ;
        RECT 47.810 -11.010 47.980 -10.840 ;
        RECT 49.420 -10.970 49.590 -10.800 ;
        RECT 52.110 -10.260 52.280 -10.090 ;
        RECT 60.530 -9.340 60.700 -9.170 ;
        RECT 61.450 -9.340 61.620 -9.170 ;
        RECT 63.080 -9.430 63.250 -9.260 ;
        RECT 70.370 -9.140 70.540 -8.970 ;
        RECT 60.020 -9.780 60.190 -9.610 ;
        RECT 54.060 -10.600 54.230 -10.430 ;
        RECT 51.010 -11.010 51.180 -10.840 ;
        RECT 52.650 -11.010 52.820 -10.840 ;
        RECT 53.560 -11.010 53.730 -10.840 ;
        RECT 55.170 -10.970 55.340 -10.800 ;
        RECT 57.860 -10.260 58.030 -10.090 ;
        RECT 66.280 -9.340 66.450 -9.170 ;
        RECT 67.200 -9.340 67.370 -9.170 ;
        RECT 68.830 -9.430 69.000 -9.260 ;
        RECT 76.120 -9.140 76.290 -8.970 ;
        RECT 65.770 -9.780 65.940 -9.610 ;
        RECT 59.810 -10.600 59.980 -10.430 ;
        RECT 56.760 -11.010 56.930 -10.840 ;
        RECT 58.400 -11.010 58.570 -10.840 ;
        RECT 59.310 -11.010 59.480 -10.840 ;
        RECT 60.920 -10.970 61.090 -10.800 ;
        RECT 63.610 -10.260 63.780 -10.090 ;
        RECT 72.030 -9.340 72.200 -9.170 ;
        RECT 72.950 -9.340 73.120 -9.170 ;
        RECT 74.580 -9.430 74.750 -9.260 ;
        RECT 81.870 -9.140 82.040 -8.970 ;
        RECT 71.520 -9.780 71.690 -9.610 ;
        RECT 65.560 -10.600 65.730 -10.430 ;
        RECT 62.510 -11.010 62.680 -10.840 ;
        RECT 64.150 -11.010 64.320 -10.840 ;
        RECT 65.060 -11.010 65.230 -10.840 ;
        RECT 66.670 -10.970 66.840 -10.800 ;
        RECT 69.360 -10.260 69.530 -10.090 ;
        RECT 77.780 -9.340 77.950 -9.170 ;
        RECT 78.700 -9.340 78.870 -9.170 ;
        RECT 80.330 -9.430 80.500 -9.260 ;
        RECT 87.620 -9.140 87.790 -8.970 ;
        RECT 77.270 -9.780 77.440 -9.610 ;
        RECT 71.310 -10.600 71.480 -10.430 ;
        RECT 68.260 -11.010 68.430 -10.840 ;
        RECT 69.900 -11.010 70.070 -10.840 ;
        RECT 70.810 -11.010 70.980 -10.840 ;
        RECT 72.420 -10.970 72.590 -10.800 ;
        RECT 75.110 -10.260 75.280 -10.090 ;
        RECT 83.530 -9.340 83.700 -9.170 ;
        RECT 84.450 -9.340 84.620 -9.170 ;
        RECT 86.080 -9.430 86.250 -9.260 ;
        RECT 93.370 -9.140 93.540 -8.970 ;
        RECT 83.020 -9.780 83.190 -9.610 ;
        RECT 77.060 -10.600 77.230 -10.430 ;
        RECT 74.010 -11.010 74.180 -10.840 ;
        RECT 75.650 -11.010 75.820 -10.840 ;
        RECT 76.560 -11.010 76.730 -10.840 ;
        RECT 78.170 -10.970 78.340 -10.800 ;
        RECT 80.860 -10.260 81.030 -10.090 ;
        RECT 89.280 -9.340 89.450 -9.170 ;
        RECT 90.200 -9.340 90.370 -9.170 ;
        RECT 91.830 -9.430 92.000 -9.260 ;
        RECT 88.770 -9.780 88.940 -9.610 ;
        RECT 82.810 -10.600 82.980 -10.430 ;
        RECT 79.760 -11.010 79.930 -10.840 ;
        RECT 81.400 -11.010 81.570 -10.840 ;
        RECT 82.310 -11.010 82.480 -10.840 ;
        RECT 83.920 -10.970 84.090 -10.800 ;
        RECT 86.610 -10.260 86.780 -10.090 ;
        RECT 88.560 -10.600 88.730 -10.430 ;
        RECT 85.510 -11.010 85.680 -10.840 ;
        RECT 87.150 -11.010 87.320 -10.840 ;
        RECT 88.060 -11.010 88.230 -10.840 ;
        RECT 89.670 -10.970 89.840 -10.800 ;
        RECT 92.360 -10.260 92.530 -10.090 ;
        RECT 94.310 -10.600 94.480 -10.430 ;
        RECT 91.260 -11.010 91.430 -10.840 ;
        RECT 92.900 -11.010 93.070 -10.840 ;
        RECT 93.810 -11.010 93.980 -10.840 ;
        RECT 3.620 -12.830 3.790 -12.660 ;
        RECT 5.310 -12.830 5.480 -12.660 ;
        RECT 6.970 -12.830 7.140 -12.660 ;
        RECT 6.010 -14.080 6.180 -13.910 ;
        RECT 9.370 -12.830 9.540 -12.660 ;
        RECT 11.060 -12.830 11.230 -12.660 ;
        RECT 12.720 -12.830 12.890 -12.660 ;
        RECT 3.410 -14.490 3.580 -14.320 ;
        RECT 3.950 -14.490 4.120 -14.320 ;
        RECT 4.080 -16.200 4.250 -16.030 ;
        RECT 5.040 -16.200 5.210 -16.030 ;
        RECT 5.570 -17.010 5.740 -16.840 ;
        RECT 11.760 -14.090 11.930 -13.920 ;
        RECT 15.120 -12.830 15.290 -12.660 ;
        RECT 16.810 -12.830 16.980 -12.660 ;
        RECT 18.470 -12.830 18.640 -12.660 ;
        RECT 6.660 -14.490 6.830 -14.320 ;
        RECT 7.200 -14.490 7.370 -14.320 ;
        RECT 9.160 -14.490 9.330 -14.320 ;
        RECT 9.700 -14.490 9.870 -14.320 ;
        RECT 6.530 -17.020 6.700 -16.850 ;
        RECT 9.830 -16.200 10.000 -16.030 ;
        RECT 10.790 -16.200 10.960 -16.030 ;
        RECT 11.320 -17.010 11.490 -16.840 ;
        RECT 17.510 -14.110 17.680 -13.940 ;
        RECT 20.870 -12.830 21.040 -12.660 ;
        RECT 22.560 -12.830 22.730 -12.660 ;
        RECT 24.220 -12.830 24.390 -12.660 ;
        RECT 12.410 -14.490 12.580 -14.320 ;
        RECT 12.950 -14.490 13.120 -14.320 ;
        RECT 14.910 -14.490 15.080 -14.320 ;
        RECT 15.450 -14.490 15.620 -14.320 ;
        RECT 12.280 -17.020 12.450 -16.850 ;
        RECT 15.580 -16.200 15.750 -16.030 ;
        RECT 16.540 -16.200 16.710 -16.030 ;
        RECT 17.070 -17.010 17.240 -16.840 ;
        RECT 23.260 -14.110 23.430 -13.940 ;
        RECT 26.620 -12.830 26.790 -12.660 ;
        RECT 28.310 -12.830 28.480 -12.660 ;
        RECT 29.970 -12.830 30.140 -12.660 ;
        RECT 18.160 -14.490 18.330 -14.320 ;
        RECT 18.700 -14.490 18.870 -14.320 ;
        RECT 20.660 -14.490 20.830 -14.320 ;
        RECT 21.200 -14.490 21.370 -14.320 ;
        RECT 18.030 -17.020 18.200 -16.850 ;
        RECT 21.330 -16.200 21.500 -16.030 ;
        RECT 22.290 -16.200 22.460 -16.030 ;
        RECT 22.820 -17.010 22.990 -16.840 ;
        RECT 29.010 -14.090 29.180 -13.920 ;
        RECT 32.370 -12.830 32.540 -12.660 ;
        RECT 34.060 -12.830 34.230 -12.660 ;
        RECT 35.720 -12.830 35.890 -12.660 ;
        RECT 23.910 -14.490 24.080 -14.320 ;
        RECT 24.450 -14.490 24.620 -14.320 ;
        RECT 26.410 -14.490 26.580 -14.320 ;
        RECT 26.950 -14.490 27.120 -14.320 ;
        RECT 23.780 -17.020 23.950 -16.850 ;
        RECT 27.080 -16.200 27.250 -16.030 ;
        RECT 28.040 -16.200 28.210 -16.030 ;
        RECT 28.570 -17.010 28.740 -16.840 ;
        RECT 34.760 -14.060 34.930 -13.890 ;
        RECT 38.120 -12.830 38.290 -12.660 ;
        RECT 39.810 -12.830 39.980 -12.660 ;
        RECT 41.470 -12.830 41.640 -12.660 ;
        RECT 29.660 -14.490 29.830 -14.320 ;
        RECT 30.200 -14.490 30.370 -14.320 ;
        RECT 32.160 -14.490 32.330 -14.320 ;
        RECT 32.700 -14.490 32.870 -14.320 ;
        RECT 29.530 -17.020 29.700 -16.850 ;
        RECT 32.830 -16.200 33.000 -16.030 ;
        RECT 33.790 -16.200 33.960 -16.030 ;
        RECT 34.320 -17.010 34.490 -16.840 ;
        RECT 40.510 -14.040 40.680 -13.870 ;
        RECT 43.870 -12.830 44.040 -12.660 ;
        RECT 45.560 -12.830 45.730 -12.660 ;
        RECT 47.220 -12.830 47.390 -12.660 ;
        RECT 35.410 -14.490 35.580 -14.320 ;
        RECT 35.950 -14.490 36.120 -14.320 ;
        RECT 37.910 -14.490 38.080 -14.320 ;
        RECT 38.450 -14.490 38.620 -14.320 ;
        RECT 35.280 -17.020 35.450 -16.850 ;
        RECT 38.580 -16.200 38.750 -16.030 ;
        RECT 39.540 -16.200 39.710 -16.030 ;
        RECT 40.070 -17.010 40.240 -16.840 ;
        RECT 46.260 -14.040 46.430 -13.870 ;
        RECT 49.620 -12.830 49.790 -12.660 ;
        RECT 51.310 -12.830 51.480 -12.660 ;
        RECT 52.970 -12.830 53.140 -12.660 ;
        RECT 41.160 -14.490 41.330 -14.320 ;
        RECT 41.700 -14.490 41.870 -14.320 ;
        RECT 43.660 -14.490 43.830 -14.320 ;
        RECT 44.200 -14.490 44.370 -14.320 ;
        RECT 41.030 -17.020 41.200 -16.850 ;
        RECT 44.330 -16.200 44.500 -16.030 ;
        RECT 45.290 -16.200 45.460 -16.030 ;
        RECT 45.820 -17.010 45.990 -16.840 ;
        RECT 52.010 -14.090 52.180 -13.920 ;
        RECT 55.370 -12.830 55.540 -12.660 ;
        RECT 57.060 -12.830 57.230 -12.660 ;
        RECT 58.720 -12.830 58.890 -12.660 ;
        RECT 46.910 -14.490 47.080 -14.320 ;
        RECT 47.450 -14.490 47.620 -14.320 ;
        RECT 49.410 -14.490 49.580 -14.320 ;
        RECT 49.950 -14.490 50.120 -14.320 ;
        RECT 46.780 -17.020 46.950 -16.850 ;
        RECT 50.080 -16.200 50.250 -16.030 ;
        RECT 51.040 -16.200 51.210 -16.030 ;
        RECT 51.570 -17.010 51.740 -16.840 ;
        RECT 57.760 -14.060 57.930 -13.890 ;
        RECT 61.120 -12.830 61.290 -12.660 ;
        RECT 62.810 -12.830 62.980 -12.660 ;
        RECT 64.470 -12.830 64.640 -12.660 ;
        RECT 52.660 -14.490 52.830 -14.320 ;
        RECT 53.200 -14.490 53.370 -14.320 ;
        RECT 55.160 -14.490 55.330 -14.320 ;
        RECT 55.700 -14.490 55.870 -14.320 ;
        RECT 52.530 -17.020 52.700 -16.850 ;
        RECT 55.830 -16.200 56.000 -16.030 ;
        RECT 56.790 -16.200 56.960 -16.030 ;
        RECT 57.320 -17.010 57.490 -16.840 ;
        RECT 63.510 -14.100 63.680 -13.930 ;
        RECT 66.870 -12.830 67.040 -12.660 ;
        RECT 68.560 -12.830 68.730 -12.660 ;
        RECT 70.220 -12.830 70.390 -12.660 ;
        RECT 58.410 -14.490 58.580 -14.320 ;
        RECT 58.950 -14.490 59.120 -14.320 ;
        RECT 60.910 -14.490 61.080 -14.320 ;
        RECT 61.450 -14.490 61.620 -14.320 ;
        RECT 58.280 -17.020 58.450 -16.850 ;
        RECT 61.580 -16.200 61.750 -16.030 ;
        RECT 62.540 -16.200 62.710 -16.030 ;
        RECT 63.070 -17.010 63.240 -16.840 ;
        RECT 69.260 -14.110 69.430 -13.940 ;
        RECT 72.620 -12.830 72.790 -12.660 ;
        RECT 74.310 -12.830 74.480 -12.660 ;
        RECT 75.970 -12.830 76.140 -12.660 ;
        RECT 64.160 -14.490 64.330 -14.320 ;
        RECT 64.700 -14.490 64.870 -14.320 ;
        RECT 66.660 -14.490 66.830 -14.320 ;
        RECT 67.200 -14.490 67.370 -14.320 ;
        RECT 64.030 -17.020 64.200 -16.850 ;
        RECT 67.330 -16.200 67.500 -16.030 ;
        RECT 68.290 -16.200 68.460 -16.030 ;
        RECT 68.820 -17.010 68.990 -16.840 ;
        RECT 75.010 -14.070 75.180 -13.900 ;
        RECT 78.370 -12.830 78.540 -12.660 ;
        RECT 80.060 -12.830 80.230 -12.660 ;
        RECT 81.720 -12.830 81.890 -12.660 ;
        RECT 69.910 -14.490 70.080 -14.320 ;
        RECT 70.450 -14.490 70.620 -14.320 ;
        RECT 72.410 -14.490 72.580 -14.320 ;
        RECT 72.950 -14.490 73.120 -14.320 ;
        RECT 69.780 -17.020 69.950 -16.850 ;
        RECT 73.080 -16.200 73.250 -16.030 ;
        RECT 74.040 -16.200 74.210 -16.030 ;
        RECT 74.570 -17.010 74.740 -16.840 ;
        RECT 80.760 -14.110 80.930 -13.940 ;
        RECT 84.120 -12.830 84.290 -12.660 ;
        RECT 85.810 -12.830 85.980 -12.660 ;
        RECT 87.470 -12.830 87.640 -12.660 ;
        RECT 75.660 -14.490 75.830 -14.320 ;
        RECT 76.200 -14.490 76.370 -14.320 ;
        RECT 78.160 -14.490 78.330 -14.320 ;
        RECT 78.700 -14.490 78.870 -14.320 ;
        RECT 75.530 -17.020 75.700 -16.850 ;
        RECT 78.830 -16.200 79.000 -16.030 ;
        RECT 79.790 -16.200 79.960 -16.030 ;
        RECT 80.320 -17.010 80.490 -16.840 ;
        RECT 86.510 -14.070 86.680 -13.900 ;
        RECT 89.870 -12.830 90.040 -12.660 ;
        RECT 91.560 -12.830 91.730 -12.660 ;
        RECT 93.220 -12.830 93.390 -12.660 ;
        RECT 81.410 -14.490 81.580 -14.320 ;
        RECT 81.950 -14.490 82.120 -14.320 ;
        RECT 83.910 -14.490 84.080 -14.320 ;
        RECT 84.450 -14.490 84.620 -14.320 ;
        RECT 81.280 -17.020 81.450 -16.850 ;
        RECT 84.580 -16.200 84.750 -16.030 ;
        RECT 85.540 -16.200 85.710 -16.030 ;
        RECT 86.070 -17.010 86.240 -16.840 ;
        RECT 92.260 -14.080 92.430 -13.910 ;
        RECT 87.160 -14.490 87.330 -14.320 ;
        RECT 87.700 -14.490 87.870 -14.320 ;
        RECT 89.660 -14.490 89.830 -14.320 ;
        RECT 90.200 -14.490 90.370 -14.320 ;
        RECT 87.030 -17.020 87.200 -16.850 ;
        RECT 90.330 -16.200 90.500 -16.030 ;
        RECT 91.290 -16.200 91.460 -16.030 ;
        RECT 91.820 -17.010 91.990 -16.840 ;
        RECT 92.910 -14.490 93.080 -14.320 ;
        RECT 93.450 -14.490 93.620 -14.320 ;
        RECT 92.780 -17.020 92.950 -16.850 ;
        RECT 3.480 -18.690 3.650 -18.520 ;
        RECT 7.160 -18.700 7.330 -18.530 ;
        RECT 9.230 -18.690 9.400 -18.520 ;
        RECT 12.910 -18.700 13.080 -18.530 ;
        RECT 14.980 -18.690 15.150 -18.520 ;
        RECT 18.660 -18.700 18.830 -18.530 ;
        RECT 20.730 -18.690 20.900 -18.520 ;
        RECT 24.410 -18.700 24.580 -18.530 ;
        RECT 26.480 -18.690 26.650 -18.520 ;
        RECT 30.160 -18.700 30.330 -18.530 ;
        RECT 32.230 -18.690 32.400 -18.520 ;
        RECT 35.910 -18.700 36.080 -18.530 ;
        RECT 37.980 -18.690 38.150 -18.520 ;
        RECT 41.660 -18.700 41.830 -18.530 ;
        RECT 43.730 -18.690 43.900 -18.520 ;
        RECT 47.410 -18.700 47.580 -18.530 ;
        RECT 49.480 -18.690 49.650 -18.520 ;
        RECT 53.160 -18.700 53.330 -18.530 ;
        RECT 55.230 -18.690 55.400 -18.520 ;
        RECT 58.910 -18.700 59.080 -18.530 ;
        RECT 60.980 -18.690 61.150 -18.520 ;
        RECT 64.660 -18.700 64.830 -18.530 ;
        RECT 66.730 -18.690 66.900 -18.520 ;
        RECT 70.410 -18.700 70.580 -18.530 ;
        RECT 72.480 -18.690 72.650 -18.520 ;
        RECT 76.160 -18.700 76.330 -18.530 ;
        RECT 78.230 -18.690 78.400 -18.520 ;
        RECT 81.910 -18.700 82.080 -18.530 ;
        RECT 83.980 -18.690 84.150 -18.520 ;
        RECT 87.660 -18.700 87.830 -18.530 ;
        RECT 89.730 -18.690 89.900 -18.520 ;
        RECT 93.410 -18.700 93.580 -18.530 ;
        RECT 8.120 -19.130 8.290 -18.960 ;
        RECT 13.870 -19.130 14.040 -18.960 ;
        RECT 19.620 -19.130 19.790 -18.960 ;
        RECT 25.370 -19.130 25.540 -18.960 ;
        RECT 31.120 -19.130 31.290 -18.960 ;
        RECT 36.870 -19.130 37.040 -18.960 ;
        RECT 42.620 -19.130 42.790 -18.960 ;
        RECT 48.370 -19.130 48.540 -18.960 ;
        RECT 54.120 -19.130 54.290 -18.960 ;
        RECT 59.870 -19.130 60.040 -18.960 ;
        RECT 65.620 -19.130 65.790 -18.960 ;
        RECT 71.370 -19.130 71.540 -18.960 ;
        RECT 77.120 -19.130 77.290 -18.960 ;
        RECT 82.870 -19.130 83.040 -18.960 ;
        RECT 88.620 -19.130 88.790 -18.960 ;
        RECT 94.230 -19.130 94.400 -18.960 ;
        RECT 4.350 -19.650 4.520 -19.480 ;
        RECT 6.230 -19.650 6.400 -19.480 ;
        RECT 10.100 -19.650 10.270 -19.480 ;
        RECT 11.980 -19.650 12.150 -19.480 ;
        RECT 15.850 -19.650 16.020 -19.480 ;
        RECT 17.730 -19.650 17.900 -19.480 ;
        RECT 21.600 -19.650 21.770 -19.480 ;
        RECT 23.480 -19.650 23.650 -19.480 ;
        RECT 27.350 -19.650 27.520 -19.480 ;
        RECT 29.230 -19.650 29.400 -19.480 ;
        RECT 33.100 -19.650 33.270 -19.480 ;
        RECT 34.980 -19.650 35.150 -19.480 ;
        RECT 38.850 -19.650 39.020 -19.480 ;
        RECT 40.730 -19.650 40.900 -19.480 ;
        RECT 44.600 -19.650 44.770 -19.480 ;
        RECT 46.480 -19.650 46.650 -19.480 ;
        RECT 50.350 -19.650 50.520 -19.480 ;
        RECT 52.230 -19.650 52.400 -19.480 ;
        RECT 56.100 -19.650 56.270 -19.480 ;
        RECT 57.980 -19.650 58.150 -19.480 ;
        RECT 61.850 -19.650 62.020 -19.480 ;
        RECT 63.730 -19.650 63.900 -19.480 ;
        RECT 67.600 -19.650 67.770 -19.480 ;
        RECT 69.480 -19.650 69.650 -19.480 ;
        RECT 73.350 -19.650 73.520 -19.480 ;
        RECT 75.230 -19.650 75.400 -19.480 ;
        RECT 79.100 -19.650 79.270 -19.480 ;
        RECT 80.980 -19.650 81.150 -19.480 ;
        RECT 84.850 -19.650 85.020 -19.480 ;
        RECT 86.730 -19.650 86.900 -19.480 ;
        RECT 90.600 -19.650 90.770 -19.480 ;
        RECT 92.480 -19.650 92.650 -19.480 ;
        RECT 4.150 -20.130 4.320 -19.960 ;
        RECT 3.140 -20.530 3.310 -20.360 ;
        RECT 5.030 -20.540 5.200 -20.370 ;
        RECT 5.550 -20.540 5.720 -20.370 ;
        RECT 6.430 -20.130 6.600 -19.960 ;
        RECT 9.900 -20.130 10.070 -19.960 ;
        RECT 3.120 -21.220 3.290 -21.050 ;
        RECT 3.640 -21.240 3.810 -21.070 ;
        RECT 5.750 -21.240 5.920 -21.070 ;
        RECT 3.140 -22.010 3.310 -21.840 ;
        RECT 7.440 -20.530 7.610 -20.360 ;
        RECT 8.890 -20.530 9.060 -20.360 ;
        RECT 10.780 -20.540 10.950 -20.370 ;
        RECT 11.300 -20.540 11.470 -20.370 ;
        RECT 12.180 -20.130 12.350 -19.960 ;
        RECT 15.650 -20.130 15.820 -19.960 ;
        RECT 7.450 -21.240 7.620 -21.070 ;
        RECT 8.870 -21.220 9.040 -21.050 ;
        RECT 9.390 -21.240 9.560 -21.070 ;
        RECT 11.500 -21.240 11.670 -21.070 ;
        RECT 7.440 -22.010 7.610 -21.840 ;
        RECT 8.890 -22.010 9.060 -21.840 ;
        RECT 13.190 -20.530 13.360 -20.360 ;
        RECT 14.640 -20.530 14.810 -20.360 ;
        RECT 16.530 -20.540 16.700 -20.370 ;
        RECT 17.050 -20.540 17.220 -20.370 ;
        RECT 17.930 -20.130 18.100 -19.960 ;
        RECT 21.400 -20.130 21.570 -19.960 ;
        RECT 13.200 -21.240 13.370 -21.070 ;
        RECT 14.620 -21.220 14.790 -21.050 ;
        RECT 15.140 -21.240 15.310 -21.070 ;
        RECT 17.250 -21.240 17.420 -21.070 ;
        RECT 13.190 -22.010 13.360 -21.840 ;
        RECT 14.640 -22.010 14.810 -21.840 ;
        RECT 18.940 -20.530 19.110 -20.360 ;
        RECT 20.390 -20.530 20.560 -20.360 ;
        RECT 22.280 -20.540 22.450 -20.370 ;
        RECT 22.800 -20.540 22.970 -20.370 ;
        RECT 23.680 -20.130 23.850 -19.960 ;
        RECT 27.150 -20.130 27.320 -19.960 ;
        RECT 18.950 -21.240 19.120 -21.070 ;
        RECT 20.370 -21.220 20.540 -21.050 ;
        RECT 20.890 -21.240 21.060 -21.070 ;
        RECT 23.000 -21.240 23.170 -21.070 ;
        RECT 18.940 -22.010 19.110 -21.840 ;
        RECT 20.390 -22.010 20.560 -21.840 ;
        RECT 24.690 -20.530 24.860 -20.360 ;
        RECT 26.140 -20.530 26.310 -20.360 ;
        RECT 28.030 -20.540 28.200 -20.370 ;
        RECT 28.550 -20.540 28.720 -20.370 ;
        RECT 29.430 -20.130 29.600 -19.960 ;
        RECT 32.900 -20.130 33.070 -19.960 ;
        RECT 24.700 -21.240 24.870 -21.070 ;
        RECT 26.120 -21.220 26.290 -21.050 ;
        RECT 26.640 -21.240 26.810 -21.070 ;
        RECT 28.750 -21.240 28.920 -21.070 ;
        RECT 24.690 -22.010 24.860 -21.840 ;
        RECT 26.140 -22.010 26.310 -21.840 ;
        RECT 30.440 -20.530 30.610 -20.360 ;
        RECT 31.890 -20.530 32.060 -20.360 ;
        RECT 33.780 -20.540 33.950 -20.370 ;
        RECT 34.300 -20.540 34.470 -20.370 ;
        RECT 35.180 -20.130 35.350 -19.960 ;
        RECT 38.650 -20.130 38.820 -19.960 ;
        RECT 30.450 -21.240 30.620 -21.070 ;
        RECT 31.870 -21.220 32.040 -21.050 ;
        RECT 32.390 -21.240 32.560 -21.070 ;
        RECT 34.500 -21.240 34.670 -21.070 ;
        RECT 30.440 -22.010 30.610 -21.840 ;
        RECT 31.890 -22.010 32.060 -21.840 ;
        RECT 36.190 -20.530 36.360 -20.360 ;
        RECT 37.640 -20.530 37.810 -20.360 ;
        RECT 39.530 -20.540 39.700 -20.370 ;
        RECT 40.050 -20.540 40.220 -20.370 ;
        RECT 40.930 -20.130 41.100 -19.960 ;
        RECT 44.400 -20.130 44.570 -19.960 ;
        RECT 36.200 -21.240 36.370 -21.070 ;
        RECT 37.620 -21.220 37.790 -21.050 ;
        RECT 38.140 -21.240 38.310 -21.070 ;
        RECT 40.250 -21.240 40.420 -21.070 ;
        RECT 36.190 -22.010 36.360 -21.840 ;
        RECT 37.640 -22.010 37.810 -21.840 ;
        RECT 41.940 -20.530 42.110 -20.360 ;
        RECT 43.390 -20.530 43.560 -20.360 ;
        RECT 45.280 -20.540 45.450 -20.370 ;
        RECT 45.800 -20.540 45.970 -20.370 ;
        RECT 46.680 -20.130 46.850 -19.960 ;
        RECT 50.150 -20.130 50.320 -19.960 ;
        RECT 41.950 -21.240 42.120 -21.070 ;
        RECT 43.370 -21.220 43.540 -21.050 ;
        RECT 43.890 -21.240 44.060 -21.070 ;
        RECT 46.000 -21.240 46.170 -21.070 ;
        RECT 41.940 -22.010 42.110 -21.840 ;
        RECT 43.390 -22.010 43.560 -21.840 ;
        RECT 47.690 -20.530 47.860 -20.360 ;
        RECT 49.140 -20.530 49.310 -20.360 ;
        RECT 51.030 -20.540 51.200 -20.370 ;
        RECT 51.550 -20.540 51.720 -20.370 ;
        RECT 52.430 -20.130 52.600 -19.960 ;
        RECT 55.900 -20.130 56.070 -19.960 ;
        RECT 47.700 -21.240 47.870 -21.070 ;
        RECT 49.120 -21.220 49.290 -21.050 ;
        RECT 49.640 -21.240 49.810 -21.070 ;
        RECT 51.750 -21.240 51.920 -21.070 ;
        RECT 47.690 -22.010 47.860 -21.840 ;
        RECT 49.140 -22.010 49.310 -21.840 ;
        RECT 53.440 -20.530 53.610 -20.360 ;
        RECT 54.890 -20.530 55.060 -20.360 ;
        RECT 56.780 -20.540 56.950 -20.370 ;
        RECT 57.300 -20.540 57.470 -20.370 ;
        RECT 58.180 -20.130 58.350 -19.960 ;
        RECT 61.650 -20.130 61.820 -19.960 ;
        RECT 53.450 -21.240 53.620 -21.070 ;
        RECT 54.870 -21.220 55.040 -21.050 ;
        RECT 55.390 -21.240 55.560 -21.070 ;
        RECT 57.500 -21.240 57.670 -21.070 ;
        RECT 53.440 -22.010 53.610 -21.840 ;
        RECT 54.890 -22.010 55.060 -21.840 ;
        RECT 59.190 -20.530 59.360 -20.360 ;
        RECT 60.640 -20.530 60.810 -20.360 ;
        RECT 62.530 -20.540 62.700 -20.370 ;
        RECT 63.050 -20.540 63.220 -20.370 ;
        RECT 63.930 -20.130 64.100 -19.960 ;
        RECT 67.400 -20.130 67.570 -19.960 ;
        RECT 59.200 -21.240 59.370 -21.070 ;
        RECT 60.620 -21.220 60.790 -21.050 ;
        RECT 61.140 -21.240 61.310 -21.070 ;
        RECT 63.250 -21.240 63.420 -21.070 ;
        RECT 59.190 -22.010 59.360 -21.840 ;
        RECT 60.640 -22.010 60.810 -21.840 ;
        RECT 64.940 -20.530 65.110 -20.360 ;
        RECT 66.390 -20.530 66.560 -20.360 ;
        RECT 68.280 -20.540 68.450 -20.370 ;
        RECT 68.800 -20.540 68.970 -20.370 ;
        RECT 69.680 -20.130 69.850 -19.960 ;
        RECT 73.150 -20.130 73.320 -19.960 ;
        RECT 64.950 -21.240 65.120 -21.070 ;
        RECT 66.370 -21.220 66.540 -21.050 ;
        RECT 66.890 -21.240 67.060 -21.070 ;
        RECT 69.000 -21.240 69.170 -21.070 ;
        RECT 64.940 -22.010 65.110 -21.840 ;
        RECT 66.390 -22.010 66.560 -21.840 ;
        RECT 70.690 -20.530 70.860 -20.360 ;
        RECT 72.140 -20.530 72.310 -20.360 ;
        RECT 74.030 -20.540 74.200 -20.370 ;
        RECT 74.550 -20.540 74.720 -20.370 ;
        RECT 75.430 -20.130 75.600 -19.960 ;
        RECT 78.900 -20.130 79.070 -19.960 ;
        RECT 70.700 -21.240 70.870 -21.070 ;
        RECT 72.120 -21.220 72.290 -21.050 ;
        RECT 72.640 -21.240 72.810 -21.070 ;
        RECT 74.750 -21.240 74.920 -21.070 ;
        RECT 70.690 -22.010 70.860 -21.840 ;
        RECT 72.140 -22.010 72.310 -21.840 ;
        RECT 76.440 -20.530 76.610 -20.360 ;
        RECT 77.890 -20.530 78.060 -20.360 ;
        RECT 79.780 -20.540 79.950 -20.370 ;
        RECT 80.300 -20.540 80.470 -20.370 ;
        RECT 81.180 -20.130 81.350 -19.960 ;
        RECT 84.650 -20.130 84.820 -19.960 ;
        RECT 76.450 -21.240 76.620 -21.070 ;
        RECT 77.870 -21.220 78.040 -21.050 ;
        RECT 78.390 -21.240 78.560 -21.070 ;
        RECT 80.500 -21.240 80.670 -21.070 ;
        RECT 76.440 -22.010 76.610 -21.840 ;
        RECT 77.890 -22.010 78.060 -21.840 ;
        RECT 82.190 -20.530 82.360 -20.360 ;
        RECT 83.640 -20.530 83.810 -20.360 ;
        RECT 85.530 -20.540 85.700 -20.370 ;
        RECT 86.050 -20.540 86.220 -20.370 ;
        RECT 86.930 -20.130 87.100 -19.960 ;
        RECT 90.400 -20.130 90.570 -19.960 ;
        RECT 82.200 -21.240 82.370 -21.070 ;
        RECT 83.620 -21.220 83.790 -21.050 ;
        RECT 84.140 -21.240 84.310 -21.070 ;
        RECT 86.250 -21.240 86.420 -21.070 ;
        RECT 82.190 -22.010 82.360 -21.840 ;
        RECT 83.640 -22.010 83.810 -21.840 ;
        RECT 87.940 -20.530 88.110 -20.360 ;
        RECT 89.390 -20.530 89.560 -20.360 ;
        RECT 91.280 -20.540 91.450 -20.370 ;
        RECT 91.800 -20.540 91.970 -20.370 ;
        RECT 92.680 -20.130 92.850 -19.960 ;
        RECT 87.950 -21.240 88.120 -21.070 ;
        RECT 89.370 -21.220 89.540 -21.050 ;
        RECT 89.890 -21.240 90.060 -21.070 ;
        RECT 92.000 -21.240 92.170 -21.070 ;
        RECT 87.940 -22.010 88.110 -21.840 ;
        RECT 89.390 -22.010 89.560 -21.840 ;
        RECT 93.690 -20.530 93.860 -20.360 ;
        RECT 93.700 -21.240 93.870 -21.070 ;
        RECT 93.690 -22.010 93.860 -21.840 ;
        RECT 6.680 -22.970 6.850 -22.800 ;
        RECT 5.290 -23.640 5.490 -23.440 ;
        RECT 9.670 -22.970 9.840 -22.800 ;
        RECT 18.190 -22.970 18.360 -22.800 ;
        RECT 7.410 -24.430 7.580 -24.260 ;
        RECT 8.960 -24.430 9.130 -24.260 ;
        RECT 21.170 -22.970 21.340 -22.800 ;
        RECT 29.690 -22.970 29.860 -22.800 ;
        RECT 32.670 -22.970 32.840 -22.800 ;
        RECT 41.190 -22.970 41.360 -22.800 ;
        RECT 44.170 -22.970 44.340 -22.800 ;
        RECT 52.690 -22.970 52.860 -22.800 ;
        RECT 30.410 -24.430 30.580 -24.260 ;
        RECT 31.950 -24.430 32.120 -24.260 ;
        RECT 55.670 -22.970 55.840 -22.800 ;
        RECT 64.190 -22.970 64.360 -22.800 ;
        RECT 41.880 -24.430 42.050 -24.260 ;
        RECT 43.470 -24.440 43.640 -24.270 ;
        RECT 67.170 -22.970 67.340 -22.800 ;
        RECT 75.690 -22.970 75.860 -22.800 ;
        RECT 53.400 -24.430 53.570 -24.260 ;
        RECT 54.950 -24.430 55.120 -24.260 ;
        RECT 78.670 -22.970 78.840 -22.800 ;
        RECT 87.190 -22.970 87.360 -22.800 ;
        RECT 64.910 -24.440 65.080 -24.270 ;
        RECT 66.440 -24.440 66.610 -24.270 ;
        RECT 90.170 -22.970 90.340 -22.800 ;
        RECT 76.420 -24.430 76.590 -24.260 ;
        RECT 77.950 -24.430 78.120 -24.260 ;
        RECT 87.910 -24.420 88.080 -24.250 ;
        RECT 89.430 -24.430 89.600 -24.260 ;
        RECT 92.090 -25.180 92.330 -24.940 ;
        RECT -37.210 -31.460 -37.040 -31.290 ;
        RECT -33.160 -31.460 -32.990 -31.290 ;
        RECT -25.710 -31.460 -25.540 -31.290 ;
        RECT -21.660 -31.460 -21.490 -31.290 ;
        RECT -13.890 -31.460 -13.720 -31.290 ;
        RECT -9.840 -31.460 -9.670 -31.290 ;
        RECT -2.080 -31.460 -1.910 -31.290 ;
        RECT 1.970 -31.460 2.140 -31.290 ;
        RECT 9.730 -31.460 9.900 -31.290 ;
        RECT 13.780 -31.460 13.950 -31.290 ;
        RECT 21.550 -31.460 21.720 -31.290 ;
        RECT 25.600 -31.460 25.770 -31.290 ;
        RECT 33.370 -31.460 33.540 -31.290 ;
        RECT 37.420 -31.460 37.590 -31.290 ;
        RECT 45.190 -31.460 45.360 -31.290 ;
        RECT 49.240 -31.460 49.410 -31.290 ;
        RECT 57.010 -31.460 57.180 -31.290 ;
        RECT 61.060 -31.460 61.230 -31.290 ;
        RECT 68.830 -31.460 69.000 -31.290 ;
        RECT 72.880 -31.460 73.050 -31.290 ;
        RECT 80.650 -31.460 80.820 -31.290 ;
        RECT 84.700 -31.460 84.870 -31.290 ;
        RECT 92.490 -31.460 92.660 -31.290 ;
        RECT 96.540 -31.460 96.710 -31.290 ;
        RECT 104.330 -31.460 104.500 -31.290 ;
        RECT 108.380 -31.460 108.550 -31.290 ;
        RECT 116.200 -31.460 116.370 -31.290 ;
        RECT 120.250 -31.460 120.420 -31.290 ;
        RECT 128.070 -31.460 128.240 -31.290 ;
        RECT 132.120 -31.460 132.290 -31.290 ;
        RECT 137.080 -31.460 137.250 -31.290 ;
        RECT 141.130 -31.460 141.300 -31.290 ;
        RECT -36.960 -33.830 -36.790 -33.660 ;
        RECT -35.170 -33.820 -35.000 -33.650 ;
        RECT -36.540 -36.060 -36.370 -35.890 ;
        RECT -33.410 -33.800 -33.240 -33.630 ;
        RECT -32.290 -33.810 -32.120 -33.640 ;
        RECT -25.460 -33.830 -25.290 -33.660 ;
        RECT -23.670 -33.820 -23.500 -33.650 ;
        RECT -24.810 -36.060 -24.640 -35.890 ;
        RECT -21.910 -33.800 -21.740 -33.630 ;
        RECT -20.790 -33.810 -20.620 -33.640 ;
        RECT -36.710 -36.500 -36.540 -36.330 ;
        RECT -37.830 -36.890 -37.660 -36.720 ;
        RECT -37.880 -37.520 -37.710 -37.350 ;
        RECT -38.230 -39.750 -38.060 -39.580 ;
        RECT -37.920 -41.550 -37.750 -41.380 ;
        RECT -37.440 -43.680 -37.270 -43.510 ;
        RECT -36.840 -39.750 -36.670 -39.580 ;
        RECT -37.830 -44.160 -37.660 -43.990 ;
        RECT -36.400 -37.490 -36.230 -37.320 ;
        RECT -36.400 -38.200 -36.230 -38.030 ;
        RECT -35.440 -38.200 -35.270 -38.030 ;
        RECT -34.910 -39.010 -34.740 -38.840 ;
        RECT -13.640 -33.830 -13.470 -33.660 ;
        RECT -11.850 -33.820 -11.680 -33.650 ;
        RECT -13.090 -36.060 -12.920 -35.890 ;
        RECT -10.090 -33.800 -9.920 -33.630 ;
        RECT -8.970 -33.810 -8.800 -33.640 ;
        RECT -33.640 -36.490 -33.470 -36.320 ;
        RECT -25.210 -36.500 -25.040 -36.330 ;
        RECT -33.950 -37.480 -33.780 -37.310 ;
        RECT -33.950 -39.020 -33.780 -38.850 ;
        RECT -32.550 -36.900 -32.380 -36.730 ;
        RECT -26.330 -36.890 -26.160 -36.720 ;
        RECT -33.510 -39.740 -33.340 -39.570 ;
        RECT -32.500 -37.510 -32.330 -37.340 ;
        RECT -26.380 -37.520 -26.210 -37.350 ;
        RECT -32.150 -39.750 -31.980 -39.580 ;
        RECT -26.730 -39.750 -26.560 -39.580 ;
        RECT -26.420 -41.550 -26.250 -41.380 ;
        RECT -25.940 -43.680 -25.770 -43.510 ;
        RECT -25.340 -39.750 -25.170 -39.580 ;
        RECT -26.330 -44.160 -26.160 -43.990 ;
        RECT -24.900 -37.490 -24.730 -37.320 ;
        RECT -24.900 -38.200 -24.730 -38.030 ;
        RECT -23.940 -38.200 -23.770 -38.030 ;
        RECT -23.410 -39.010 -23.240 -38.840 ;
        RECT -1.830 -33.830 -1.660 -33.660 ;
        RECT -0.040 -33.820 0.130 -33.650 ;
        RECT -1.280 -36.060 -1.110 -35.890 ;
        RECT 1.720 -33.800 1.890 -33.630 ;
        RECT 2.840 -33.810 3.010 -33.640 ;
        RECT -22.140 -36.490 -21.970 -36.320 ;
        RECT -13.390 -36.500 -13.220 -36.330 ;
        RECT -22.450 -37.480 -22.280 -37.310 ;
        RECT -22.450 -39.020 -22.280 -38.850 ;
        RECT -21.050 -36.900 -20.880 -36.730 ;
        RECT -14.510 -36.890 -14.340 -36.720 ;
        RECT -22.010 -39.740 -21.840 -39.570 ;
        RECT -21.000 -37.510 -20.830 -37.340 ;
        RECT -14.560 -37.520 -14.390 -37.350 ;
        RECT -20.650 -39.750 -20.480 -39.580 ;
        RECT -14.910 -39.750 -14.740 -39.580 ;
        RECT -14.600 -41.550 -14.430 -41.380 ;
        RECT -14.120 -43.680 -13.950 -43.510 ;
        RECT -13.520 -39.750 -13.350 -39.580 ;
        RECT -14.510 -44.160 -14.340 -43.990 ;
        RECT -13.080 -37.490 -12.910 -37.320 ;
        RECT -13.080 -38.200 -12.910 -38.030 ;
        RECT -12.120 -38.200 -11.950 -38.030 ;
        RECT -11.590 -39.010 -11.420 -38.840 ;
        RECT 9.980 -33.830 10.150 -33.660 ;
        RECT 11.770 -33.820 11.940 -33.650 ;
        RECT 10.580 -36.060 10.750 -35.890 ;
        RECT 13.530 -33.800 13.700 -33.630 ;
        RECT 14.650 -33.810 14.820 -33.640 ;
        RECT -10.320 -36.490 -10.150 -36.320 ;
        RECT -1.580 -36.500 -1.410 -36.330 ;
        RECT -10.630 -37.480 -10.460 -37.310 ;
        RECT -10.630 -39.020 -10.460 -38.850 ;
        RECT -9.230 -36.900 -9.060 -36.730 ;
        RECT -2.700 -36.890 -2.530 -36.720 ;
        RECT -10.190 -39.740 -10.020 -39.570 ;
        RECT -9.180 -37.510 -9.010 -37.340 ;
        RECT -2.750 -37.520 -2.580 -37.350 ;
        RECT -8.830 -39.750 -8.660 -39.580 ;
        RECT -3.100 -39.750 -2.930 -39.580 ;
        RECT -2.790 -41.550 -2.620 -41.380 ;
        RECT -2.310 -43.680 -2.140 -43.510 ;
        RECT -1.710 -39.750 -1.540 -39.580 ;
        RECT -2.700 -44.160 -2.530 -43.990 ;
        RECT -1.270 -37.490 -1.100 -37.320 ;
        RECT -1.270 -38.200 -1.100 -38.030 ;
        RECT -0.310 -38.200 -0.140 -38.030 ;
        RECT 0.220 -39.010 0.390 -38.840 ;
        RECT 21.800 -33.830 21.970 -33.660 ;
        RECT 23.590 -33.820 23.760 -33.650 ;
        RECT 22.420 -36.060 22.590 -35.890 ;
        RECT 25.350 -33.800 25.520 -33.630 ;
        RECT 26.470 -33.810 26.640 -33.640 ;
        RECT 1.490 -36.490 1.660 -36.320 ;
        RECT 10.230 -36.500 10.400 -36.330 ;
        RECT 1.180 -37.480 1.350 -37.310 ;
        RECT 1.180 -39.020 1.350 -38.850 ;
        RECT 2.580 -36.900 2.750 -36.730 ;
        RECT 9.110 -36.890 9.280 -36.720 ;
        RECT 1.620 -39.740 1.790 -39.570 ;
        RECT 2.630 -37.510 2.800 -37.340 ;
        RECT 9.060 -37.520 9.230 -37.350 ;
        RECT 2.980 -39.750 3.150 -39.580 ;
        RECT 8.710 -39.750 8.880 -39.580 ;
        RECT 9.020 -41.550 9.190 -41.380 ;
        RECT 9.500 -43.680 9.670 -43.510 ;
        RECT 10.100 -39.750 10.270 -39.580 ;
        RECT 9.110 -44.160 9.280 -43.990 ;
        RECT 10.540 -37.490 10.710 -37.320 ;
        RECT 10.540 -38.200 10.710 -38.030 ;
        RECT 11.500 -38.200 11.670 -38.030 ;
        RECT 12.030 -39.010 12.200 -38.840 ;
        RECT 33.620 -33.830 33.790 -33.660 ;
        RECT 35.410 -33.820 35.580 -33.650 ;
        RECT 34.100 -36.060 34.270 -35.890 ;
        RECT 37.170 -33.800 37.340 -33.630 ;
        RECT 38.290 -33.810 38.460 -33.640 ;
        RECT 13.300 -36.490 13.470 -36.320 ;
        RECT 22.050 -36.500 22.220 -36.330 ;
        RECT 12.990 -37.480 13.160 -37.310 ;
        RECT 12.990 -39.020 13.160 -38.850 ;
        RECT 14.390 -36.900 14.560 -36.730 ;
        RECT 20.930 -36.890 21.100 -36.720 ;
        RECT 13.430 -39.740 13.600 -39.570 ;
        RECT 14.440 -37.510 14.610 -37.340 ;
        RECT 20.880 -37.520 21.050 -37.350 ;
        RECT 14.790 -39.750 14.960 -39.580 ;
        RECT 20.530 -39.750 20.700 -39.580 ;
        RECT 20.840 -41.550 21.010 -41.380 ;
        RECT 21.320 -43.680 21.490 -43.510 ;
        RECT 21.920 -39.750 22.090 -39.580 ;
        RECT 20.930 -44.160 21.100 -43.990 ;
        RECT 22.360 -37.490 22.530 -37.320 ;
        RECT 22.360 -38.200 22.530 -38.030 ;
        RECT 23.320 -38.200 23.490 -38.030 ;
        RECT 23.850 -39.010 24.020 -38.840 ;
        RECT 45.440 -33.830 45.610 -33.660 ;
        RECT 47.230 -33.820 47.400 -33.650 ;
        RECT 45.990 -36.060 46.160 -35.890 ;
        RECT 48.990 -33.800 49.160 -33.630 ;
        RECT 50.110 -33.810 50.280 -33.640 ;
        RECT 25.120 -36.490 25.290 -36.320 ;
        RECT 33.870 -36.500 34.040 -36.330 ;
        RECT 24.810 -37.480 24.980 -37.310 ;
        RECT 24.810 -39.020 24.980 -38.850 ;
        RECT 26.210 -36.900 26.380 -36.730 ;
        RECT 32.750 -36.890 32.920 -36.720 ;
        RECT 25.250 -39.740 25.420 -39.570 ;
        RECT 26.260 -37.510 26.430 -37.340 ;
        RECT 32.700 -37.520 32.870 -37.350 ;
        RECT 26.610 -39.750 26.780 -39.580 ;
        RECT 32.350 -39.750 32.520 -39.580 ;
        RECT 32.660 -41.550 32.830 -41.380 ;
        RECT 33.140 -43.680 33.310 -43.510 ;
        RECT 33.740 -39.750 33.910 -39.580 ;
        RECT 32.750 -44.160 32.920 -43.990 ;
        RECT 34.180 -37.490 34.350 -37.320 ;
        RECT 34.180 -38.200 34.350 -38.030 ;
        RECT 35.140 -38.200 35.310 -38.030 ;
        RECT 35.670 -39.010 35.840 -38.840 ;
        RECT 57.260 -33.830 57.430 -33.660 ;
        RECT 59.050 -33.820 59.220 -33.650 ;
        RECT 57.770 -36.060 57.940 -35.890 ;
        RECT 60.810 -33.800 60.980 -33.630 ;
        RECT 61.930 -33.810 62.100 -33.640 ;
        RECT 36.940 -36.490 37.110 -36.320 ;
        RECT 45.690 -36.500 45.860 -36.330 ;
        RECT 36.630 -37.480 36.800 -37.310 ;
        RECT 36.630 -39.020 36.800 -38.850 ;
        RECT 38.030 -36.900 38.200 -36.730 ;
        RECT 44.570 -36.890 44.740 -36.720 ;
        RECT 37.070 -39.740 37.240 -39.570 ;
        RECT 38.080 -37.510 38.250 -37.340 ;
        RECT 44.520 -37.520 44.690 -37.350 ;
        RECT 38.430 -39.750 38.600 -39.580 ;
        RECT 44.170 -39.750 44.340 -39.580 ;
        RECT 44.480 -41.550 44.650 -41.380 ;
        RECT 44.960 -43.680 45.130 -43.510 ;
        RECT 45.560 -39.750 45.730 -39.580 ;
        RECT 44.570 -44.160 44.740 -43.990 ;
        RECT 46.000 -37.490 46.170 -37.320 ;
        RECT 46.000 -38.200 46.170 -38.030 ;
        RECT 46.960 -38.200 47.130 -38.030 ;
        RECT 47.490 -39.010 47.660 -38.840 ;
        RECT 69.080 -33.830 69.250 -33.660 ;
        RECT 70.870 -33.820 71.040 -33.650 ;
        RECT 69.660 -36.060 69.830 -35.890 ;
        RECT 72.630 -33.800 72.800 -33.630 ;
        RECT 73.750 -33.810 73.920 -33.640 ;
        RECT 48.760 -36.490 48.930 -36.320 ;
        RECT 57.510 -36.500 57.680 -36.330 ;
        RECT 48.450 -37.480 48.620 -37.310 ;
        RECT 48.450 -39.020 48.620 -38.850 ;
        RECT 49.850 -36.900 50.020 -36.730 ;
        RECT 56.390 -36.890 56.560 -36.720 ;
        RECT 48.890 -39.740 49.060 -39.570 ;
        RECT 49.900 -37.510 50.070 -37.340 ;
        RECT 56.340 -37.520 56.510 -37.350 ;
        RECT 50.250 -39.750 50.420 -39.580 ;
        RECT 55.990 -39.750 56.160 -39.580 ;
        RECT 56.300 -41.550 56.470 -41.380 ;
        RECT 56.780 -43.680 56.950 -43.510 ;
        RECT 57.380 -39.750 57.550 -39.580 ;
        RECT 56.390 -44.160 56.560 -43.990 ;
        RECT 57.820 -37.490 57.990 -37.320 ;
        RECT 57.820 -38.200 57.990 -38.030 ;
        RECT 58.780 -38.200 58.950 -38.030 ;
        RECT 59.310 -39.010 59.480 -38.840 ;
        RECT 80.900 -33.830 81.070 -33.660 ;
        RECT 82.690 -33.820 82.860 -33.650 ;
        RECT 81.320 -36.060 81.490 -35.890 ;
        RECT 84.450 -33.800 84.620 -33.630 ;
        RECT 85.570 -33.810 85.740 -33.640 ;
        RECT 60.580 -36.490 60.750 -36.320 ;
        RECT 69.330 -36.500 69.500 -36.330 ;
        RECT 60.270 -37.480 60.440 -37.310 ;
        RECT 60.270 -39.020 60.440 -38.850 ;
        RECT 61.670 -36.900 61.840 -36.730 ;
        RECT 68.210 -36.890 68.380 -36.720 ;
        RECT 60.710 -39.740 60.880 -39.570 ;
        RECT 61.720 -37.510 61.890 -37.340 ;
        RECT 68.160 -37.520 68.330 -37.350 ;
        RECT 62.070 -39.750 62.240 -39.580 ;
        RECT 67.810 -39.750 67.980 -39.580 ;
        RECT 68.120 -41.550 68.290 -41.380 ;
        RECT 68.600 -43.680 68.770 -43.510 ;
        RECT 69.200 -39.750 69.370 -39.580 ;
        RECT 68.210 -44.160 68.380 -43.990 ;
        RECT 69.640 -37.490 69.810 -37.320 ;
        RECT 69.640 -38.200 69.810 -38.030 ;
        RECT 70.600 -38.200 70.770 -38.030 ;
        RECT 71.130 -39.010 71.300 -38.840 ;
        RECT 92.740 -33.830 92.910 -33.660 ;
        RECT 94.530 -33.820 94.700 -33.650 ;
        RECT 93.340 -36.060 93.510 -35.890 ;
        RECT 96.290 -33.800 96.460 -33.630 ;
        RECT 97.410 -33.810 97.580 -33.640 ;
        RECT 72.400 -36.490 72.570 -36.320 ;
        RECT 81.150 -36.500 81.320 -36.330 ;
        RECT 72.090 -37.480 72.260 -37.310 ;
        RECT 72.090 -39.020 72.260 -38.850 ;
        RECT 73.490 -36.900 73.660 -36.730 ;
        RECT 80.030 -36.890 80.200 -36.720 ;
        RECT 72.530 -39.740 72.700 -39.570 ;
        RECT 73.540 -37.510 73.710 -37.340 ;
        RECT 79.980 -37.520 80.150 -37.350 ;
        RECT 73.890 -39.750 74.060 -39.580 ;
        RECT 79.630 -39.750 79.800 -39.580 ;
        RECT 79.940 -41.550 80.110 -41.380 ;
        RECT 80.420 -43.680 80.590 -43.510 ;
        RECT 81.020 -39.750 81.190 -39.580 ;
        RECT 80.030 -44.160 80.200 -43.990 ;
        RECT 81.460 -37.490 81.630 -37.320 ;
        RECT 81.460 -38.200 81.630 -38.030 ;
        RECT 82.420 -38.200 82.590 -38.030 ;
        RECT 82.950 -39.010 83.120 -38.840 ;
        RECT 104.580 -33.830 104.750 -33.660 ;
        RECT 106.370 -33.820 106.540 -33.650 ;
        RECT 105.070 -36.060 105.240 -35.890 ;
        RECT 108.130 -33.800 108.300 -33.630 ;
        RECT 109.250 -33.810 109.420 -33.640 ;
        RECT 84.220 -36.490 84.390 -36.320 ;
        RECT 92.990 -36.500 93.160 -36.330 ;
        RECT 83.910 -37.480 84.080 -37.310 ;
        RECT 83.910 -39.020 84.080 -38.850 ;
        RECT 85.310 -36.900 85.480 -36.730 ;
        RECT 91.870 -36.890 92.040 -36.720 ;
        RECT 84.350 -39.740 84.520 -39.570 ;
        RECT 85.360 -37.510 85.530 -37.340 ;
        RECT 91.820 -37.520 91.990 -37.350 ;
        RECT 85.710 -39.750 85.880 -39.580 ;
        RECT 91.470 -39.750 91.640 -39.580 ;
        RECT 91.780 -41.550 91.950 -41.380 ;
        RECT 92.260 -43.680 92.430 -43.510 ;
        RECT 92.860 -39.750 93.030 -39.580 ;
        RECT 91.870 -44.160 92.040 -43.990 ;
        RECT 93.300 -37.490 93.470 -37.320 ;
        RECT 93.300 -38.200 93.470 -38.030 ;
        RECT 94.260 -38.200 94.430 -38.030 ;
        RECT 94.790 -39.010 94.960 -38.840 ;
        RECT 116.450 -33.830 116.620 -33.660 ;
        RECT 118.240 -33.820 118.410 -33.650 ;
        RECT 116.790 -36.060 116.960 -35.890 ;
        RECT 120.000 -33.800 120.170 -33.630 ;
        RECT 121.120 -33.810 121.290 -33.640 ;
        RECT 96.060 -36.490 96.230 -36.320 ;
        RECT 104.830 -36.500 105.000 -36.330 ;
        RECT 95.750 -37.480 95.920 -37.310 ;
        RECT 95.750 -39.020 95.920 -38.850 ;
        RECT 97.150 -36.900 97.320 -36.730 ;
        RECT 103.710 -36.890 103.880 -36.720 ;
        RECT 96.190 -39.740 96.360 -39.570 ;
        RECT 97.200 -37.510 97.370 -37.340 ;
        RECT 103.660 -37.520 103.830 -37.350 ;
        RECT 97.550 -39.750 97.720 -39.580 ;
        RECT 103.310 -39.750 103.480 -39.580 ;
        RECT 103.620 -41.550 103.790 -41.380 ;
        RECT 104.100 -43.680 104.270 -43.510 ;
        RECT 104.700 -39.750 104.870 -39.580 ;
        RECT 103.710 -44.160 103.880 -43.990 ;
        RECT 105.140 -37.490 105.310 -37.320 ;
        RECT 105.140 -38.200 105.310 -38.030 ;
        RECT 106.100 -38.200 106.270 -38.030 ;
        RECT 106.630 -39.010 106.800 -38.840 ;
        RECT 128.320 -33.830 128.490 -33.660 ;
        RECT 130.110 -33.820 130.280 -33.650 ;
        RECT 128.950 -36.060 129.120 -35.890 ;
        RECT 131.870 -33.800 132.040 -33.630 ;
        RECT 132.990 -33.810 133.160 -33.640 ;
        RECT 107.900 -36.490 108.070 -36.320 ;
        RECT 116.700 -36.500 116.870 -36.330 ;
        RECT 107.590 -37.480 107.760 -37.310 ;
        RECT 107.590 -39.020 107.760 -38.850 ;
        RECT 108.990 -36.900 109.160 -36.730 ;
        RECT 115.580 -36.890 115.750 -36.720 ;
        RECT 108.030 -39.740 108.200 -39.570 ;
        RECT 109.040 -37.510 109.210 -37.340 ;
        RECT 115.530 -37.520 115.700 -37.350 ;
        RECT 109.390 -39.750 109.560 -39.580 ;
        RECT 115.180 -39.750 115.350 -39.580 ;
        RECT 115.490 -41.550 115.660 -41.380 ;
        RECT 115.970 -43.680 116.140 -43.510 ;
        RECT 116.570 -39.750 116.740 -39.580 ;
        RECT 115.580 -44.160 115.750 -43.990 ;
        RECT 117.010 -37.490 117.180 -37.320 ;
        RECT 117.010 -38.200 117.180 -38.030 ;
        RECT 117.970 -38.200 118.140 -38.030 ;
        RECT 118.500 -39.010 118.670 -38.840 ;
        RECT 137.330 -33.830 137.500 -33.660 ;
        RECT 139.120 -33.820 139.290 -33.650 ;
        RECT 137.970 -36.060 138.140 -35.890 ;
        RECT 140.880 -33.800 141.050 -33.630 ;
        RECT 142.000 -33.810 142.170 -33.640 ;
        RECT 119.770 -36.490 119.940 -36.320 ;
        RECT 128.570 -36.500 128.740 -36.330 ;
        RECT 119.460 -37.480 119.630 -37.310 ;
        RECT 119.460 -39.020 119.630 -38.850 ;
        RECT 120.860 -36.900 121.030 -36.730 ;
        RECT 127.450 -36.890 127.620 -36.720 ;
        RECT 119.900 -39.740 120.070 -39.570 ;
        RECT 120.910 -37.510 121.080 -37.340 ;
        RECT 127.400 -37.520 127.570 -37.350 ;
        RECT 121.260 -39.750 121.430 -39.580 ;
        RECT 127.050 -39.750 127.220 -39.580 ;
        RECT 127.360 -41.550 127.530 -41.380 ;
        RECT 127.840 -43.680 128.010 -43.510 ;
        RECT 128.440 -39.750 128.610 -39.580 ;
        RECT 127.450 -44.160 127.620 -43.990 ;
        RECT 128.880 -37.490 129.050 -37.320 ;
        RECT 128.880 -38.200 129.050 -38.030 ;
        RECT 129.840 -38.200 130.010 -38.030 ;
        RECT 130.370 -39.010 130.540 -38.840 ;
        RECT 131.640 -36.490 131.810 -36.320 ;
        RECT 137.580 -36.500 137.750 -36.330 ;
        RECT 131.330 -37.480 131.500 -37.310 ;
        RECT 131.330 -39.020 131.500 -38.850 ;
        RECT 132.730 -36.900 132.900 -36.730 ;
        RECT 136.460 -36.890 136.630 -36.720 ;
        RECT 131.770 -39.740 131.940 -39.570 ;
        RECT 132.780 -37.510 132.950 -37.340 ;
        RECT 136.410 -37.520 136.580 -37.350 ;
        RECT 133.130 -39.750 133.300 -39.580 ;
        RECT 136.060 -39.750 136.230 -39.580 ;
        RECT 136.370 -41.550 136.540 -41.380 ;
        RECT 136.850 -43.680 137.020 -43.510 ;
        RECT 137.450 -39.750 137.620 -39.580 ;
        RECT 136.460 -44.160 136.630 -43.990 ;
        RECT 137.890 -37.490 138.060 -37.320 ;
        RECT 137.890 -38.200 138.060 -38.030 ;
        RECT 138.850 -38.200 139.020 -38.030 ;
        RECT 139.380 -39.010 139.550 -38.840 ;
        RECT 140.650 -36.490 140.820 -36.320 ;
        RECT 140.340 -37.480 140.510 -37.310 ;
        RECT 140.340 -39.020 140.510 -38.850 ;
        RECT 141.740 -36.900 141.910 -36.730 ;
        RECT 140.780 -39.740 140.950 -39.570 ;
        RECT 141.790 -37.510 141.960 -37.340 ;
        RECT 142.140 -39.750 142.310 -39.580 ;
        RECT -32.820 -45.170 -32.650 -45.000 ;
        RECT -21.320 -45.170 -21.150 -45.000 ;
        RECT -9.500 -45.170 -9.330 -45.000 ;
        RECT 2.310 -45.170 2.480 -45.000 ;
        RECT 14.120 -45.170 14.290 -45.000 ;
        RECT 25.940 -45.170 26.110 -45.000 ;
        RECT 37.760 -45.170 37.930 -45.000 ;
        RECT 49.580 -45.170 49.750 -45.000 ;
        RECT 61.400 -45.170 61.570 -45.000 ;
        RECT 73.220 -45.170 73.390 -45.000 ;
        RECT 85.040 -45.170 85.210 -45.000 ;
        RECT 96.880 -45.170 97.050 -45.000 ;
        RECT 108.720 -45.170 108.890 -45.000 ;
        RECT 120.590 -45.170 120.760 -45.000 ;
        RECT 132.460 -45.170 132.630 -45.000 ;
        RECT 141.470 -45.170 141.640 -45.000 ;
        RECT -37.440 -46.570 -37.270 -46.400 ;
        RECT -37.830 -48.710 -37.660 -48.540 ;
        RECT -38.230 -50.500 -38.060 -50.330 ;
        RECT -37.880 -52.730 -37.710 -52.560 ;
        RECT -36.840 -50.500 -36.670 -50.330 ;
        RECT -37.830 -53.360 -37.660 -53.190 ;
        RECT -36.400 -52.050 -36.230 -51.880 ;
        RECT -36.400 -52.760 -36.230 -52.590 ;
        RECT -36.710 -53.750 -36.540 -53.580 ;
        RECT -35.440 -52.050 -35.270 -51.880 ;
        RECT -34.910 -51.240 -34.740 -51.070 ;
        RECT -36.320 -54.180 -36.150 -54.010 ;
        RECT -33.950 -51.230 -33.780 -51.060 ;
        RECT -33.950 -52.770 -33.780 -52.600 ;
        RECT -32.150 -45.570 -31.980 -45.400 ;
        RECT -25.940 -46.570 -25.770 -46.400 ;
        RECT -26.330 -48.710 -26.160 -48.540 ;
        RECT -33.510 -50.510 -33.340 -50.340 ;
        RECT -32.150 -50.500 -31.980 -50.330 ;
        RECT -26.730 -50.500 -26.560 -50.330 ;
        RECT -32.500 -52.740 -32.330 -52.570 ;
        RECT -26.380 -52.730 -26.210 -52.560 ;
        RECT -25.340 -50.500 -25.170 -50.330 ;
        RECT -32.550 -53.350 -32.380 -53.180 ;
        RECT -26.330 -53.360 -26.160 -53.190 ;
        RECT -24.900 -52.050 -24.730 -51.880 ;
        RECT -24.900 -52.760 -24.730 -52.590 ;
        RECT -33.640 -53.760 -33.470 -53.590 ;
        RECT -25.210 -53.750 -25.040 -53.580 ;
        RECT -23.940 -52.050 -23.770 -51.880 ;
        RECT -23.410 -51.240 -23.240 -51.070 ;
        RECT -22.450 -51.230 -22.280 -51.060 ;
        RECT -22.450 -52.770 -22.280 -52.600 ;
        RECT -20.650 -45.560 -20.480 -45.390 ;
        RECT -14.120 -46.570 -13.950 -46.400 ;
        RECT -14.510 -48.710 -14.340 -48.540 ;
        RECT -22.010 -50.510 -21.840 -50.340 ;
        RECT -20.650 -50.500 -20.480 -50.330 ;
        RECT -14.910 -50.500 -14.740 -50.330 ;
        RECT -21.000 -52.740 -20.830 -52.570 ;
        RECT -14.560 -52.730 -14.390 -52.560 ;
        RECT -13.520 -50.500 -13.350 -50.330 ;
        RECT -21.050 -53.350 -20.880 -53.180 ;
        RECT -14.510 -53.360 -14.340 -53.190 ;
        RECT -13.080 -52.050 -12.910 -51.880 ;
        RECT -13.080 -52.760 -12.910 -52.590 ;
        RECT -22.140 -53.760 -21.970 -53.590 ;
        RECT -13.390 -53.750 -13.220 -53.580 ;
        RECT -12.120 -52.050 -11.950 -51.880 ;
        RECT -11.590 -51.240 -11.420 -51.070 ;
        RECT -36.960 -56.420 -36.790 -56.250 ;
        RECT -35.170 -56.430 -35.000 -56.260 ;
        RECT -33.410 -56.450 -33.240 -56.280 ;
        RECT -25.010 -54.190 -24.840 -54.020 ;
        RECT -10.630 -51.230 -10.460 -51.060 ;
        RECT -10.630 -52.770 -10.460 -52.600 ;
        RECT -8.830 -45.590 -8.660 -45.420 ;
        RECT -2.310 -46.570 -2.140 -46.400 ;
        RECT -2.700 -48.710 -2.530 -48.540 ;
        RECT -10.190 -50.510 -10.020 -50.340 ;
        RECT -8.830 -50.500 -8.660 -50.330 ;
        RECT -3.100 -50.500 -2.930 -50.330 ;
        RECT -9.180 -52.740 -9.010 -52.570 ;
        RECT -2.750 -52.730 -2.580 -52.560 ;
        RECT -1.710 -50.500 -1.540 -50.330 ;
        RECT -9.230 -53.350 -9.060 -53.180 ;
        RECT -2.700 -53.360 -2.530 -53.190 ;
        RECT -1.270 -52.050 -1.100 -51.880 ;
        RECT -1.270 -52.760 -1.100 -52.590 ;
        RECT -10.320 -53.760 -10.150 -53.590 ;
        RECT -1.580 -53.750 -1.410 -53.580 ;
        RECT -0.310 -52.050 -0.140 -51.880 ;
        RECT 0.220 -51.240 0.390 -51.070 ;
        RECT -32.290 -56.430 -32.120 -56.260 ;
        RECT -25.460 -56.420 -25.290 -56.250 ;
        RECT -23.670 -56.430 -23.500 -56.260 ;
        RECT -21.910 -56.450 -21.740 -56.280 ;
        RECT -13.200 -54.190 -13.030 -54.020 ;
        RECT 1.180 -51.230 1.350 -51.060 ;
        RECT 1.180 -52.770 1.350 -52.600 ;
        RECT 2.980 -45.560 3.150 -45.390 ;
        RECT 9.500 -46.570 9.670 -46.400 ;
        RECT 9.110 -48.710 9.280 -48.540 ;
        RECT 1.620 -50.510 1.790 -50.340 ;
        RECT 2.980 -50.500 3.150 -50.330 ;
        RECT 8.710 -50.500 8.880 -50.330 ;
        RECT 2.630 -52.740 2.800 -52.570 ;
        RECT 9.060 -52.730 9.230 -52.560 ;
        RECT 10.100 -50.500 10.270 -50.330 ;
        RECT 2.580 -53.350 2.750 -53.180 ;
        RECT 9.110 -53.360 9.280 -53.190 ;
        RECT 10.540 -52.050 10.710 -51.880 ;
        RECT 10.540 -52.760 10.710 -52.590 ;
        RECT 1.490 -53.760 1.660 -53.590 ;
        RECT 10.230 -53.750 10.400 -53.580 ;
        RECT 11.500 -52.050 11.670 -51.880 ;
        RECT 12.030 -51.240 12.200 -51.070 ;
        RECT -20.790 -56.430 -20.620 -56.260 ;
        RECT -13.640 -56.420 -13.470 -56.250 ;
        RECT -11.850 -56.430 -11.680 -56.260 ;
        RECT -10.090 -56.450 -9.920 -56.280 ;
        RECT -1.480 -54.190 -1.310 -54.020 ;
        RECT 12.990 -51.230 13.160 -51.060 ;
        RECT 12.990 -52.770 13.160 -52.600 ;
        RECT 14.790 -45.560 14.960 -45.390 ;
        RECT 21.320 -46.570 21.490 -46.400 ;
        RECT 20.930 -48.710 21.100 -48.540 ;
        RECT 13.430 -50.510 13.600 -50.340 ;
        RECT 14.790 -50.500 14.960 -50.330 ;
        RECT 20.530 -50.500 20.700 -50.330 ;
        RECT 14.440 -52.740 14.610 -52.570 ;
        RECT 20.880 -52.730 21.050 -52.560 ;
        RECT 21.920 -50.500 22.090 -50.330 ;
        RECT 14.390 -53.350 14.560 -53.180 ;
        RECT 20.930 -53.360 21.100 -53.190 ;
        RECT 22.360 -52.050 22.530 -51.880 ;
        RECT 22.360 -52.760 22.530 -52.590 ;
        RECT 13.300 -53.760 13.470 -53.590 ;
        RECT 22.050 -53.750 22.220 -53.580 ;
        RECT 23.320 -52.050 23.490 -51.880 ;
        RECT 23.850 -51.240 24.020 -51.070 ;
        RECT -8.970 -56.430 -8.800 -56.260 ;
        RECT -1.830 -56.420 -1.660 -56.250 ;
        RECT -0.040 -56.430 0.130 -56.260 ;
        RECT 1.720 -56.450 1.890 -56.280 ;
        RECT 10.300 -54.190 10.470 -54.020 ;
        RECT 24.810 -51.230 24.980 -51.060 ;
        RECT 24.810 -52.770 24.980 -52.600 ;
        RECT 26.610 -45.560 26.780 -45.390 ;
        RECT 33.140 -46.570 33.310 -46.400 ;
        RECT 32.750 -48.710 32.920 -48.540 ;
        RECT 25.250 -50.510 25.420 -50.340 ;
        RECT 26.610 -50.500 26.780 -50.330 ;
        RECT 32.350 -50.500 32.520 -50.330 ;
        RECT 26.260 -52.740 26.430 -52.570 ;
        RECT 32.700 -52.730 32.870 -52.560 ;
        RECT 33.740 -50.500 33.910 -50.330 ;
        RECT 26.210 -53.350 26.380 -53.180 ;
        RECT 32.750 -53.360 32.920 -53.190 ;
        RECT 34.180 -52.050 34.350 -51.880 ;
        RECT 34.180 -52.760 34.350 -52.590 ;
        RECT 25.120 -53.760 25.290 -53.590 ;
        RECT 33.870 -53.750 34.040 -53.580 ;
        RECT 35.140 -52.050 35.310 -51.880 ;
        RECT 35.670 -51.240 35.840 -51.070 ;
        RECT 2.840 -56.430 3.010 -56.260 ;
        RECT 9.980 -56.420 10.150 -56.250 ;
        RECT 11.770 -56.430 11.940 -56.260 ;
        RECT 13.530 -56.450 13.700 -56.280 ;
        RECT 22.180 -54.190 22.350 -54.020 ;
        RECT 36.630 -51.230 36.800 -51.060 ;
        RECT 36.630 -52.770 36.800 -52.600 ;
        RECT 38.430 -45.560 38.600 -45.390 ;
        RECT 44.960 -46.570 45.130 -46.400 ;
        RECT 44.570 -48.710 44.740 -48.540 ;
        RECT 37.070 -50.510 37.240 -50.340 ;
        RECT 38.430 -50.500 38.600 -50.330 ;
        RECT 44.170 -50.500 44.340 -50.330 ;
        RECT 38.080 -52.740 38.250 -52.570 ;
        RECT 44.520 -52.730 44.690 -52.560 ;
        RECT 45.560 -50.500 45.730 -50.330 ;
        RECT 38.030 -53.350 38.200 -53.180 ;
        RECT 44.570 -53.360 44.740 -53.190 ;
        RECT 46.000 -52.050 46.170 -51.880 ;
        RECT 46.000 -52.760 46.170 -52.590 ;
        RECT 36.940 -53.760 37.110 -53.590 ;
        RECT 45.690 -53.750 45.860 -53.580 ;
        RECT 46.960 -52.050 47.130 -51.880 ;
        RECT 47.490 -51.240 47.660 -51.070 ;
        RECT 14.650 -56.430 14.820 -56.260 ;
        RECT 21.800 -56.420 21.970 -56.250 ;
        RECT 23.590 -56.430 23.760 -56.260 ;
        RECT 25.350 -56.450 25.520 -56.280 ;
        RECT 34.090 -54.190 34.260 -54.020 ;
        RECT 48.450 -51.230 48.620 -51.060 ;
        RECT 48.450 -52.770 48.620 -52.600 ;
        RECT 50.250 -45.560 50.420 -45.390 ;
        RECT 56.780 -46.570 56.950 -46.400 ;
        RECT 56.390 -48.710 56.560 -48.540 ;
        RECT 48.890 -50.510 49.060 -50.340 ;
        RECT 50.250 -50.500 50.420 -50.330 ;
        RECT 55.990 -50.500 56.160 -50.330 ;
        RECT 49.900 -52.740 50.070 -52.570 ;
        RECT 56.340 -52.730 56.510 -52.560 ;
        RECT 57.380 -50.500 57.550 -50.330 ;
        RECT 49.850 -53.350 50.020 -53.180 ;
        RECT 56.390 -53.360 56.560 -53.190 ;
        RECT 57.820 -52.050 57.990 -51.880 ;
        RECT 57.820 -52.760 57.990 -52.590 ;
        RECT 48.760 -53.760 48.930 -53.590 ;
        RECT 57.510 -53.750 57.680 -53.580 ;
        RECT 58.780 -52.050 58.950 -51.880 ;
        RECT 59.310 -51.240 59.480 -51.070 ;
        RECT 26.470 -56.430 26.640 -56.260 ;
        RECT 33.620 -56.420 33.790 -56.250 ;
        RECT 35.410 -56.430 35.580 -56.260 ;
        RECT 37.170 -56.450 37.340 -56.280 ;
        RECT 45.910 -54.190 46.080 -54.020 ;
        RECT 60.270 -51.230 60.440 -51.060 ;
        RECT 60.270 -52.770 60.440 -52.600 ;
        RECT 62.070 -45.560 62.240 -45.390 ;
        RECT 68.600 -46.570 68.770 -46.400 ;
        RECT 68.210 -48.710 68.380 -48.540 ;
        RECT 60.710 -50.510 60.880 -50.340 ;
        RECT 62.070 -50.500 62.240 -50.330 ;
        RECT 67.810 -50.500 67.980 -50.330 ;
        RECT 61.720 -52.740 61.890 -52.570 ;
        RECT 68.160 -52.730 68.330 -52.560 ;
        RECT 69.200 -50.500 69.370 -50.330 ;
        RECT 61.670 -53.350 61.840 -53.180 ;
        RECT 68.210 -53.360 68.380 -53.190 ;
        RECT 69.640 -52.050 69.810 -51.880 ;
        RECT 69.640 -52.760 69.810 -52.590 ;
        RECT 60.580 -53.760 60.750 -53.590 ;
        RECT 69.330 -53.750 69.500 -53.580 ;
        RECT 70.600 -52.050 70.770 -51.880 ;
        RECT 71.130 -51.240 71.300 -51.070 ;
        RECT 38.290 -56.430 38.460 -56.260 ;
        RECT 45.440 -56.420 45.610 -56.250 ;
        RECT 47.230 -56.430 47.400 -56.260 ;
        RECT 48.990 -56.450 49.160 -56.280 ;
        RECT 57.600 -54.190 57.770 -54.020 ;
        RECT 72.090 -51.230 72.260 -51.060 ;
        RECT 72.090 -52.770 72.260 -52.600 ;
        RECT 73.890 -45.560 74.060 -45.390 ;
        RECT 80.420 -46.570 80.590 -46.400 ;
        RECT 80.030 -48.710 80.200 -48.540 ;
        RECT 72.530 -50.510 72.700 -50.340 ;
        RECT 73.890 -50.500 74.060 -50.330 ;
        RECT 79.630 -50.500 79.800 -50.330 ;
        RECT 73.540 -52.740 73.710 -52.570 ;
        RECT 79.980 -52.730 80.150 -52.560 ;
        RECT 81.020 -50.500 81.190 -50.330 ;
        RECT 73.490 -53.350 73.660 -53.180 ;
        RECT 80.030 -53.360 80.200 -53.190 ;
        RECT 81.460 -52.050 81.630 -51.880 ;
        RECT 81.460 -52.760 81.630 -52.590 ;
        RECT 72.400 -53.760 72.570 -53.590 ;
        RECT 81.150 -53.750 81.320 -53.580 ;
        RECT 82.420 -52.050 82.590 -51.880 ;
        RECT 82.950 -51.240 83.120 -51.070 ;
        RECT 50.110 -56.430 50.280 -56.260 ;
        RECT 57.260 -56.420 57.430 -56.250 ;
        RECT 59.050 -56.430 59.220 -56.260 ;
        RECT 60.810 -56.450 60.980 -56.280 ;
        RECT 69.480 -54.190 69.650 -54.020 ;
        RECT 83.910 -51.230 84.080 -51.060 ;
        RECT 83.910 -52.770 84.080 -52.600 ;
        RECT 85.710 -45.560 85.880 -45.390 ;
        RECT 92.260 -46.570 92.430 -46.400 ;
        RECT 91.870 -48.710 92.040 -48.540 ;
        RECT 84.350 -50.510 84.520 -50.340 ;
        RECT 85.710 -50.500 85.880 -50.330 ;
        RECT 91.470 -50.500 91.640 -50.330 ;
        RECT 85.360 -52.740 85.530 -52.570 ;
        RECT 91.820 -52.730 91.990 -52.560 ;
        RECT 92.860 -50.500 93.030 -50.330 ;
        RECT 85.310 -53.350 85.480 -53.180 ;
        RECT 91.870 -53.360 92.040 -53.190 ;
        RECT 93.300 -52.050 93.470 -51.880 ;
        RECT 93.300 -52.760 93.470 -52.590 ;
        RECT 84.220 -53.760 84.390 -53.590 ;
        RECT 92.990 -53.750 93.160 -53.580 ;
        RECT 94.260 -52.050 94.430 -51.880 ;
        RECT 94.790 -51.240 94.960 -51.070 ;
        RECT 61.930 -56.430 62.100 -56.260 ;
        RECT 69.080 -56.420 69.250 -56.250 ;
        RECT 70.870 -56.430 71.040 -56.260 ;
        RECT 72.630 -56.450 72.800 -56.280 ;
        RECT 81.270 -54.190 81.440 -54.020 ;
        RECT 95.750 -51.230 95.920 -51.060 ;
        RECT 95.750 -52.770 95.920 -52.600 ;
        RECT 97.550 -45.560 97.720 -45.390 ;
        RECT 104.100 -46.570 104.270 -46.400 ;
        RECT 103.710 -48.710 103.880 -48.540 ;
        RECT 96.190 -50.510 96.360 -50.340 ;
        RECT 97.550 -50.500 97.720 -50.330 ;
        RECT 103.310 -50.500 103.480 -50.330 ;
        RECT 97.200 -52.740 97.370 -52.570 ;
        RECT 103.660 -52.730 103.830 -52.560 ;
        RECT 104.700 -50.500 104.870 -50.330 ;
        RECT 97.150 -53.350 97.320 -53.180 ;
        RECT 103.710 -53.360 103.880 -53.190 ;
        RECT 105.140 -52.050 105.310 -51.880 ;
        RECT 105.140 -52.760 105.310 -52.590 ;
        RECT 96.060 -53.760 96.230 -53.590 ;
        RECT 104.830 -53.750 105.000 -53.580 ;
        RECT 106.100 -52.050 106.270 -51.880 ;
        RECT 106.630 -51.240 106.800 -51.070 ;
        RECT 73.750 -56.430 73.920 -56.260 ;
        RECT 80.900 -56.420 81.070 -56.250 ;
        RECT 82.690 -56.430 82.860 -56.260 ;
        RECT 84.450 -56.450 84.620 -56.280 ;
        RECT 93.150 -54.190 93.320 -54.020 ;
        RECT 107.590 -51.230 107.760 -51.060 ;
        RECT 107.590 -52.770 107.760 -52.600 ;
        RECT 109.390 -45.570 109.560 -45.400 ;
        RECT 115.970 -46.570 116.140 -46.400 ;
        RECT 115.580 -48.710 115.750 -48.540 ;
        RECT 108.030 -50.510 108.200 -50.340 ;
        RECT 109.390 -50.500 109.560 -50.330 ;
        RECT 115.180 -50.500 115.350 -50.330 ;
        RECT 109.040 -52.740 109.210 -52.570 ;
        RECT 115.530 -52.730 115.700 -52.560 ;
        RECT 116.570 -50.500 116.740 -50.330 ;
        RECT 108.990 -53.350 109.160 -53.180 ;
        RECT 115.580 -53.360 115.750 -53.190 ;
        RECT 117.010 -52.050 117.180 -51.880 ;
        RECT 117.010 -52.760 117.180 -52.590 ;
        RECT 107.900 -53.760 108.070 -53.590 ;
        RECT 116.700 -53.750 116.870 -53.580 ;
        RECT 117.970 -52.050 118.140 -51.880 ;
        RECT 118.500 -51.240 118.670 -51.070 ;
        RECT 85.570 -56.430 85.740 -56.260 ;
        RECT 92.740 -56.420 92.910 -56.250 ;
        RECT 94.530 -56.430 94.700 -56.260 ;
        RECT 96.290 -56.450 96.460 -56.280 ;
        RECT 104.920 -54.190 105.090 -54.020 ;
        RECT 119.460 -51.230 119.630 -51.060 ;
        RECT 119.460 -52.770 119.630 -52.600 ;
        RECT 121.260 -45.560 121.430 -45.390 ;
        RECT 127.840 -46.570 128.010 -46.400 ;
        RECT 127.450 -48.710 127.620 -48.540 ;
        RECT 119.900 -50.510 120.070 -50.340 ;
        RECT 121.260 -50.500 121.430 -50.330 ;
        RECT 127.050 -50.500 127.220 -50.330 ;
        RECT 120.910 -52.740 121.080 -52.570 ;
        RECT 127.400 -52.730 127.570 -52.560 ;
        RECT 128.440 -50.500 128.610 -50.330 ;
        RECT 120.860 -53.350 121.030 -53.180 ;
        RECT 127.450 -53.360 127.620 -53.190 ;
        RECT 128.880 -52.050 129.050 -51.880 ;
        RECT 128.880 -52.760 129.050 -52.590 ;
        RECT 119.770 -53.760 119.940 -53.590 ;
        RECT 128.570 -53.750 128.740 -53.580 ;
        RECT 129.840 -52.050 130.010 -51.880 ;
        RECT 130.370 -51.240 130.540 -51.070 ;
        RECT 97.410 -56.430 97.580 -56.260 ;
        RECT 104.580 -56.420 104.750 -56.250 ;
        RECT 106.370 -56.430 106.540 -56.260 ;
        RECT 108.130 -56.450 108.300 -56.280 ;
        RECT 116.700 -54.190 116.870 -54.020 ;
        RECT 131.330 -51.230 131.500 -51.060 ;
        RECT 131.330 -52.770 131.500 -52.600 ;
        RECT 133.130 -45.560 133.300 -45.390 ;
        RECT 136.850 -46.570 137.020 -46.400 ;
        RECT 136.460 -48.710 136.630 -48.540 ;
        RECT 131.770 -50.510 131.940 -50.340 ;
        RECT 133.130 -50.500 133.300 -50.330 ;
        RECT 136.060 -50.500 136.230 -50.330 ;
        RECT 132.780 -52.740 132.950 -52.570 ;
        RECT 136.410 -52.730 136.580 -52.560 ;
        RECT 137.450 -50.500 137.620 -50.330 ;
        RECT 132.730 -53.350 132.900 -53.180 ;
        RECT 136.460 -53.360 136.630 -53.190 ;
        RECT 137.890 -52.050 138.060 -51.880 ;
        RECT 137.890 -52.760 138.060 -52.590 ;
        RECT 131.640 -53.760 131.810 -53.590 ;
        RECT 137.580 -53.750 137.750 -53.580 ;
        RECT 138.850 -52.050 139.020 -51.880 ;
        RECT 139.380 -51.240 139.550 -51.070 ;
        RECT 109.250 -56.430 109.420 -56.260 ;
        RECT 116.450 -56.420 116.620 -56.250 ;
        RECT 118.240 -56.430 118.410 -56.260 ;
        RECT 120.000 -56.450 120.170 -56.280 ;
        RECT 128.510 -54.190 128.680 -54.020 ;
        RECT 140.340 -51.230 140.510 -51.060 ;
        RECT 140.340 -52.770 140.510 -52.600 ;
        RECT 142.140 -45.560 142.310 -45.390 ;
        RECT 140.780 -50.510 140.950 -50.340 ;
        RECT 142.140 -50.500 142.310 -50.330 ;
        RECT 141.790 -52.740 141.960 -52.570 ;
        RECT 141.740 -53.350 141.910 -53.180 ;
        RECT 140.650 -53.760 140.820 -53.590 ;
        RECT 121.120 -56.430 121.290 -56.260 ;
        RECT 128.320 -56.420 128.490 -56.250 ;
        RECT 130.110 -56.430 130.280 -56.260 ;
        RECT 131.870 -56.450 132.040 -56.280 ;
        RECT 137.780 -54.190 137.950 -54.020 ;
        RECT 132.990 -56.430 133.160 -56.260 ;
        RECT 137.330 -56.420 137.500 -56.250 ;
        RECT 139.120 -56.430 139.290 -56.260 ;
        RECT 140.880 -56.450 141.050 -56.280 ;
        RECT 142.000 -56.430 142.170 -56.260 ;
        RECT -37.210 -58.790 -37.040 -58.620 ;
        RECT -33.160 -58.790 -32.990 -58.620 ;
        RECT -25.710 -58.790 -25.540 -58.620 ;
        RECT -21.660 -58.790 -21.490 -58.620 ;
        RECT -13.890 -58.790 -13.720 -58.620 ;
        RECT -9.840 -58.790 -9.670 -58.620 ;
        RECT -2.080 -58.790 -1.910 -58.620 ;
        RECT 1.970 -58.790 2.140 -58.620 ;
        RECT 9.730 -58.790 9.900 -58.620 ;
        RECT 13.780 -58.790 13.950 -58.620 ;
        RECT 21.550 -58.790 21.720 -58.620 ;
        RECT 25.600 -58.790 25.770 -58.620 ;
        RECT 33.370 -58.790 33.540 -58.620 ;
        RECT 37.420 -58.790 37.590 -58.620 ;
        RECT 45.190 -58.790 45.360 -58.620 ;
        RECT 49.240 -58.790 49.410 -58.620 ;
        RECT 57.010 -58.790 57.180 -58.620 ;
        RECT 61.060 -58.790 61.230 -58.620 ;
        RECT 68.830 -58.790 69.000 -58.620 ;
        RECT 72.880 -58.790 73.050 -58.620 ;
        RECT 80.650 -58.790 80.820 -58.620 ;
        RECT 84.700 -58.790 84.870 -58.620 ;
        RECT 92.490 -58.790 92.660 -58.620 ;
        RECT 96.540 -58.790 96.710 -58.620 ;
        RECT 104.330 -58.790 104.500 -58.620 ;
        RECT 108.380 -58.790 108.550 -58.620 ;
        RECT 116.200 -58.790 116.370 -58.620 ;
        RECT 120.250 -58.790 120.420 -58.620 ;
        RECT 128.070 -58.790 128.240 -58.620 ;
        RECT 132.120 -58.790 132.290 -58.620 ;
        RECT 137.080 -58.790 137.250 -58.620 ;
        RECT 141.130 -58.790 141.300 -58.620 ;
        RECT -36.960 -61.160 -36.790 -60.990 ;
        RECT -35.170 -61.150 -35.000 -60.980 ;
        RECT -36.340 -63.390 -36.170 -63.220 ;
        RECT -33.410 -61.130 -33.240 -60.960 ;
        RECT -32.300 -61.140 -32.130 -60.970 ;
        RECT -25.460 -61.160 -25.290 -60.990 ;
        RECT -23.670 -61.150 -23.500 -60.980 ;
        RECT -24.860 -63.390 -24.690 -63.220 ;
        RECT -21.910 -61.130 -21.740 -60.960 ;
        RECT -20.800 -61.140 -20.630 -60.970 ;
        RECT -36.710 -63.830 -36.540 -63.660 ;
        RECT -37.830 -64.220 -37.660 -64.050 ;
        RECT -37.880 -64.850 -37.710 -64.680 ;
        RECT -37.830 -66.280 -37.660 -66.110 ;
        RECT -38.230 -67.080 -38.060 -66.910 ;
        RECT -37.840 -68.870 -37.670 -68.700 ;
        RECT -37.440 -71.010 -37.270 -70.840 ;
        RECT -36.840 -67.080 -36.670 -66.910 ;
        RECT -36.400 -64.820 -36.230 -64.650 ;
        RECT -36.400 -65.530 -36.230 -65.360 ;
        RECT -35.440 -65.530 -35.270 -65.360 ;
        RECT -34.910 -66.340 -34.740 -66.170 ;
        RECT -13.640 -61.160 -13.470 -60.990 ;
        RECT -11.850 -61.150 -11.680 -60.980 ;
        RECT -13.050 -63.390 -12.880 -63.220 ;
        RECT -10.090 -61.130 -9.920 -60.960 ;
        RECT -8.980 -61.140 -8.810 -60.970 ;
        RECT -33.640 -63.820 -33.470 -63.650 ;
        RECT -25.210 -63.830 -25.040 -63.660 ;
        RECT -33.950 -64.810 -33.780 -64.640 ;
        RECT -33.950 -66.350 -33.780 -66.180 ;
        RECT -32.550 -64.230 -32.380 -64.060 ;
        RECT -26.330 -64.220 -26.160 -64.050 ;
        RECT -33.510 -67.070 -33.340 -66.900 ;
        RECT -32.500 -64.840 -32.330 -64.670 ;
        RECT -26.380 -64.850 -26.210 -64.680 ;
        RECT -26.330 -66.280 -26.160 -66.110 ;
        RECT -32.150 -67.080 -31.980 -66.910 ;
        RECT -26.730 -67.080 -26.560 -66.910 ;
        RECT -26.340 -68.870 -26.170 -68.700 ;
        RECT -25.940 -71.010 -25.770 -70.840 ;
        RECT -25.340 -67.080 -25.170 -66.910 ;
        RECT -24.900 -64.820 -24.730 -64.650 ;
        RECT -24.900 -65.530 -24.730 -65.360 ;
        RECT -23.940 -65.530 -23.770 -65.360 ;
        RECT -23.410 -66.340 -23.240 -66.170 ;
        RECT -1.830 -61.160 -1.660 -60.990 ;
        RECT -0.040 -61.150 0.130 -60.980 ;
        RECT -1.300 -63.390 -1.130 -63.220 ;
        RECT 1.720 -61.130 1.890 -60.960 ;
        RECT 2.830 -61.140 3.000 -60.970 ;
        RECT -22.140 -63.820 -21.970 -63.650 ;
        RECT -13.390 -63.830 -13.220 -63.660 ;
        RECT -22.450 -64.810 -22.280 -64.640 ;
        RECT -22.450 -66.350 -22.280 -66.180 ;
        RECT -21.050 -64.230 -20.880 -64.060 ;
        RECT -14.510 -64.220 -14.340 -64.050 ;
        RECT -22.010 -67.070 -21.840 -66.900 ;
        RECT -21.000 -64.840 -20.830 -64.670 ;
        RECT -14.560 -64.850 -14.390 -64.680 ;
        RECT -14.510 -66.280 -14.340 -66.110 ;
        RECT -20.650 -67.080 -20.480 -66.910 ;
        RECT -14.910 -67.080 -14.740 -66.910 ;
        RECT -14.520 -68.870 -14.350 -68.700 ;
        RECT -14.120 -71.010 -13.950 -70.840 ;
        RECT -13.520 -67.080 -13.350 -66.910 ;
        RECT -13.080 -64.820 -12.910 -64.650 ;
        RECT -13.080 -65.530 -12.910 -65.360 ;
        RECT -12.120 -65.530 -11.950 -65.360 ;
        RECT -11.590 -66.340 -11.420 -66.170 ;
        RECT 9.980 -61.160 10.150 -60.990 ;
        RECT 11.770 -61.150 11.940 -60.980 ;
        RECT 10.580 -63.390 10.750 -63.220 ;
        RECT 13.530 -61.130 13.700 -60.960 ;
        RECT 14.640 -61.140 14.810 -60.970 ;
        RECT -10.320 -63.820 -10.150 -63.650 ;
        RECT -1.580 -63.830 -1.410 -63.660 ;
        RECT -10.630 -64.810 -10.460 -64.640 ;
        RECT -10.630 -66.350 -10.460 -66.180 ;
        RECT -9.230 -64.230 -9.060 -64.060 ;
        RECT -2.700 -64.220 -2.530 -64.050 ;
        RECT -10.190 -67.070 -10.020 -66.900 ;
        RECT -9.180 -64.840 -9.010 -64.670 ;
        RECT -2.750 -64.850 -2.580 -64.680 ;
        RECT -2.700 -66.280 -2.530 -66.110 ;
        RECT -8.830 -67.080 -8.660 -66.910 ;
        RECT -3.100 -67.080 -2.930 -66.910 ;
        RECT -2.710 -68.870 -2.540 -68.700 ;
        RECT -2.310 -71.010 -2.140 -70.840 ;
        RECT -1.710 -67.080 -1.540 -66.910 ;
        RECT -1.270 -64.820 -1.100 -64.650 ;
        RECT -1.270 -65.530 -1.100 -65.360 ;
        RECT -0.310 -65.530 -0.140 -65.360 ;
        RECT 0.220 -66.340 0.390 -66.170 ;
        RECT 21.800 -61.160 21.970 -60.990 ;
        RECT 23.590 -61.150 23.760 -60.980 ;
        RECT 22.420 -63.390 22.590 -63.220 ;
        RECT 25.350 -61.130 25.520 -60.960 ;
        RECT 26.460 -61.140 26.630 -60.970 ;
        RECT 1.490 -63.820 1.660 -63.650 ;
        RECT 10.230 -63.830 10.400 -63.660 ;
        RECT 1.180 -64.810 1.350 -64.640 ;
        RECT 1.180 -66.350 1.350 -66.180 ;
        RECT 2.580 -64.230 2.750 -64.060 ;
        RECT 9.110 -64.220 9.280 -64.050 ;
        RECT 1.620 -67.070 1.790 -66.900 ;
        RECT 2.630 -64.840 2.800 -64.670 ;
        RECT 9.060 -64.850 9.230 -64.680 ;
        RECT 9.110 -66.280 9.280 -66.110 ;
        RECT 2.980 -67.080 3.150 -66.910 ;
        RECT 8.710 -67.080 8.880 -66.910 ;
        RECT 9.100 -68.870 9.270 -68.700 ;
        RECT 9.500 -71.010 9.670 -70.840 ;
        RECT 10.100 -67.080 10.270 -66.910 ;
        RECT 10.540 -64.820 10.710 -64.650 ;
        RECT 10.540 -65.530 10.710 -65.360 ;
        RECT 11.500 -65.530 11.670 -65.360 ;
        RECT 12.030 -66.340 12.200 -66.170 ;
        RECT 33.620 -61.160 33.790 -60.990 ;
        RECT 35.410 -61.150 35.580 -60.980 ;
        RECT 34.130 -63.390 34.300 -63.220 ;
        RECT 37.170 -61.130 37.340 -60.960 ;
        RECT 38.280 -61.140 38.450 -60.970 ;
        RECT 13.300 -63.820 13.470 -63.650 ;
        RECT 22.050 -63.830 22.220 -63.660 ;
        RECT 12.990 -64.810 13.160 -64.640 ;
        RECT 12.990 -66.350 13.160 -66.180 ;
        RECT 14.390 -64.230 14.560 -64.060 ;
        RECT 20.930 -64.220 21.100 -64.050 ;
        RECT 13.430 -67.070 13.600 -66.900 ;
        RECT 14.440 -64.840 14.610 -64.670 ;
        RECT 20.880 -64.850 21.050 -64.680 ;
        RECT 20.930 -66.280 21.100 -66.110 ;
        RECT 14.790 -67.080 14.960 -66.910 ;
        RECT 20.530 -67.080 20.700 -66.910 ;
        RECT 20.920 -68.870 21.090 -68.700 ;
        RECT 21.320 -71.010 21.490 -70.840 ;
        RECT 21.920 -67.080 22.090 -66.910 ;
        RECT 22.360 -64.820 22.530 -64.650 ;
        RECT 22.360 -65.530 22.530 -65.360 ;
        RECT 23.320 -65.530 23.490 -65.360 ;
        RECT 23.850 -66.340 24.020 -66.170 ;
        RECT 45.440 -61.160 45.610 -60.990 ;
        RECT 47.230 -61.150 47.400 -60.980 ;
        RECT 46.000 -63.390 46.170 -63.220 ;
        RECT 48.990 -61.130 49.160 -60.960 ;
        RECT 50.100 -61.140 50.270 -60.970 ;
        RECT 25.120 -63.820 25.290 -63.650 ;
        RECT 33.870 -63.830 34.040 -63.660 ;
        RECT 24.810 -64.810 24.980 -64.640 ;
        RECT 24.810 -66.350 24.980 -66.180 ;
        RECT 26.210 -64.230 26.380 -64.060 ;
        RECT 32.750 -64.220 32.920 -64.050 ;
        RECT 25.250 -67.070 25.420 -66.900 ;
        RECT 26.260 -64.840 26.430 -64.670 ;
        RECT 32.700 -64.850 32.870 -64.680 ;
        RECT 32.750 -66.280 32.920 -66.110 ;
        RECT 26.610 -67.080 26.780 -66.910 ;
        RECT 32.350 -67.080 32.520 -66.910 ;
        RECT 32.740 -68.870 32.910 -68.700 ;
        RECT 33.140 -71.010 33.310 -70.840 ;
        RECT 33.740 -67.080 33.910 -66.910 ;
        RECT 34.180 -64.820 34.350 -64.650 ;
        RECT 34.180 -65.530 34.350 -65.360 ;
        RECT 35.140 -65.530 35.310 -65.360 ;
        RECT 35.670 -66.340 35.840 -66.170 ;
        RECT 57.260 -61.160 57.430 -60.990 ;
        RECT 59.050 -61.150 59.220 -60.980 ;
        RECT 57.880 -63.390 58.050 -63.220 ;
        RECT 60.810 -61.130 60.980 -60.960 ;
        RECT 61.920 -61.140 62.090 -60.970 ;
        RECT 36.940 -63.820 37.110 -63.650 ;
        RECT 45.690 -63.830 45.860 -63.660 ;
        RECT 36.630 -64.810 36.800 -64.640 ;
        RECT 36.630 -66.350 36.800 -66.180 ;
        RECT 38.030 -64.230 38.200 -64.060 ;
        RECT 44.570 -64.220 44.740 -64.050 ;
        RECT 37.070 -67.070 37.240 -66.900 ;
        RECT 38.080 -64.840 38.250 -64.670 ;
        RECT 44.520 -64.850 44.690 -64.680 ;
        RECT 44.570 -66.280 44.740 -66.110 ;
        RECT 38.430 -67.080 38.600 -66.910 ;
        RECT 44.170 -67.080 44.340 -66.910 ;
        RECT 44.560 -68.870 44.730 -68.700 ;
        RECT 44.960 -71.010 45.130 -70.840 ;
        RECT 45.560 -67.080 45.730 -66.910 ;
        RECT 46.000 -64.820 46.170 -64.650 ;
        RECT 46.000 -65.530 46.170 -65.360 ;
        RECT 46.960 -65.530 47.130 -65.360 ;
        RECT 47.490 -66.340 47.660 -66.170 ;
        RECT 69.080 -61.160 69.250 -60.990 ;
        RECT 70.870 -61.150 71.040 -60.980 ;
        RECT 69.550 -63.390 69.720 -63.220 ;
        RECT 72.630 -61.130 72.800 -60.960 ;
        RECT 73.740 -61.140 73.910 -60.970 ;
        RECT 48.760 -63.820 48.930 -63.650 ;
        RECT 57.510 -63.830 57.680 -63.660 ;
        RECT 48.450 -64.810 48.620 -64.640 ;
        RECT 48.450 -66.350 48.620 -66.180 ;
        RECT 49.850 -64.230 50.020 -64.060 ;
        RECT 56.390 -64.220 56.560 -64.050 ;
        RECT 48.890 -67.070 49.060 -66.900 ;
        RECT 49.900 -64.840 50.070 -64.670 ;
        RECT 56.340 -64.850 56.510 -64.680 ;
        RECT 56.390 -66.280 56.560 -66.110 ;
        RECT 50.250 -67.080 50.420 -66.910 ;
        RECT 55.990 -67.080 56.160 -66.910 ;
        RECT 56.380 -68.870 56.550 -68.700 ;
        RECT 56.780 -71.010 56.950 -70.840 ;
        RECT 57.380 -67.080 57.550 -66.910 ;
        RECT 57.820 -64.820 57.990 -64.650 ;
        RECT 57.820 -65.530 57.990 -65.360 ;
        RECT 58.780 -65.530 58.950 -65.360 ;
        RECT 59.310 -66.340 59.480 -66.170 ;
        RECT 80.900 -61.160 81.070 -60.990 ;
        RECT 82.690 -61.150 82.860 -60.980 ;
        RECT 81.370 -63.390 81.540 -63.220 ;
        RECT 84.450 -61.130 84.620 -60.960 ;
        RECT 85.560 -61.140 85.730 -60.970 ;
        RECT 60.580 -63.820 60.750 -63.650 ;
        RECT 69.330 -63.830 69.500 -63.660 ;
        RECT 60.270 -64.810 60.440 -64.640 ;
        RECT 60.270 -66.350 60.440 -66.180 ;
        RECT 61.670 -64.230 61.840 -64.060 ;
        RECT 68.210 -64.220 68.380 -64.050 ;
        RECT 60.710 -67.070 60.880 -66.900 ;
        RECT 61.720 -64.840 61.890 -64.670 ;
        RECT 68.160 -64.850 68.330 -64.680 ;
        RECT 68.210 -66.280 68.380 -66.110 ;
        RECT 62.070 -67.080 62.240 -66.910 ;
        RECT 67.810 -67.080 67.980 -66.910 ;
        RECT 68.200 -68.870 68.370 -68.700 ;
        RECT 68.600 -71.010 68.770 -70.840 ;
        RECT 69.200 -67.080 69.370 -66.910 ;
        RECT 69.640 -64.820 69.810 -64.650 ;
        RECT 69.640 -65.530 69.810 -65.360 ;
        RECT 70.600 -65.530 70.770 -65.360 ;
        RECT 71.130 -66.340 71.300 -66.170 ;
        RECT 92.740 -61.160 92.910 -60.990 ;
        RECT 94.530 -61.150 94.700 -60.980 ;
        RECT 93.230 -63.390 93.400 -63.220 ;
        RECT 96.290 -61.130 96.460 -60.960 ;
        RECT 97.400 -61.140 97.570 -60.970 ;
        RECT 72.400 -63.820 72.570 -63.650 ;
        RECT 81.150 -63.830 81.320 -63.660 ;
        RECT 72.090 -64.810 72.260 -64.640 ;
        RECT 72.090 -66.350 72.260 -66.180 ;
        RECT 73.490 -64.230 73.660 -64.060 ;
        RECT 80.030 -64.220 80.200 -64.050 ;
        RECT 72.530 -67.070 72.700 -66.900 ;
        RECT 73.540 -64.840 73.710 -64.670 ;
        RECT 79.980 -64.850 80.150 -64.680 ;
        RECT 80.030 -66.280 80.200 -66.110 ;
        RECT 73.890 -67.080 74.060 -66.910 ;
        RECT 79.630 -67.080 79.800 -66.910 ;
        RECT 80.020 -68.870 80.190 -68.700 ;
        RECT 80.420 -71.010 80.590 -70.840 ;
        RECT 81.020 -67.080 81.190 -66.910 ;
        RECT 81.460 -64.820 81.630 -64.650 ;
        RECT 81.460 -65.530 81.630 -65.360 ;
        RECT 82.420 -65.530 82.590 -65.360 ;
        RECT 82.950 -66.340 83.120 -66.170 ;
        RECT 104.580 -61.160 104.750 -60.990 ;
        RECT 106.370 -61.150 106.540 -60.980 ;
        RECT 104.990 -63.390 105.160 -63.220 ;
        RECT 108.130 -61.130 108.300 -60.960 ;
        RECT 109.240 -61.140 109.410 -60.970 ;
        RECT 84.220 -63.820 84.390 -63.650 ;
        RECT 92.990 -63.830 93.160 -63.660 ;
        RECT 83.910 -64.810 84.080 -64.640 ;
        RECT 83.910 -66.350 84.080 -66.180 ;
        RECT 85.310 -64.230 85.480 -64.060 ;
        RECT 91.870 -64.220 92.040 -64.050 ;
        RECT 84.350 -67.070 84.520 -66.900 ;
        RECT 85.360 -64.840 85.530 -64.670 ;
        RECT 91.820 -64.850 91.990 -64.680 ;
        RECT 91.870 -66.280 92.040 -66.110 ;
        RECT 85.710 -67.080 85.880 -66.910 ;
        RECT 91.470 -67.080 91.640 -66.910 ;
        RECT 91.860 -68.870 92.030 -68.700 ;
        RECT 92.260 -71.010 92.430 -70.840 ;
        RECT 92.860 -67.080 93.030 -66.910 ;
        RECT 93.300 -64.820 93.470 -64.650 ;
        RECT 93.300 -65.530 93.470 -65.360 ;
        RECT 94.260 -65.530 94.430 -65.360 ;
        RECT 94.790 -66.340 94.960 -66.170 ;
        RECT 116.450 -61.160 116.620 -60.990 ;
        RECT 118.240 -61.150 118.410 -60.980 ;
        RECT 116.780 -63.390 116.950 -63.220 ;
        RECT 120.000 -61.130 120.170 -60.960 ;
        RECT 121.110 -61.140 121.280 -60.970 ;
        RECT 96.060 -63.820 96.230 -63.650 ;
        RECT 104.830 -63.830 105.000 -63.660 ;
        RECT 95.750 -64.810 95.920 -64.640 ;
        RECT 95.750 -66.350 95.920 -66.180 ;
        RECT 97.150 -64.230 97.320 -64.060 ;
        RECT 103.710 -64.220 103.880 -64.050 ;
        RECT 96.190 -67.070 96.360 -66.900 ;
        RECT 97.200 -64.840 97.370 -64.670 ;
        RECT 103.660 -64.850 103.830 -64.680 ;
        RECT 103.710 -66.280 103.880 -66.110 ;
        RECT 97.550 -67.080 97.720 -66.910 ;
        RECT 103.310 -67.080 103.480 -66.910 ;
        RECT 103.700 -68.870 103.870 -68.700 ;
        RECT 104.100 -71.010 104.270 -70.840 ;
        RECT 104.700 -67.080 104.870 -66.910 ;
        RECT 105.140 -64.820 105.310 -64.650 ;
        RECT 105.140 -65.530 105.310 -65.360 ;
        RECT 106.100 -65.530 106.270 -65.360 ;
        RECT 106.630 -66.340 106.800 -66.170 ;
        RECT 128.320 -61.160 128.490 -60.990 ;
        RECT 130.110 -61.150 130.280 -60.980 ;
        RECT 128.800 -63.390 128.970 -63.220 ;
        RECT 131.870 -61.130 132.040 -60.960 ;
        RECT 132.980 -61.140 133.150 -60.970 ;
        RECT 107.900 -63.820 108.070 -63.650 ;
        RECT 116.700 -63.830 116.870 -63.660 ;
        RECT 107.590 -64.810 107.760 -64.640 ;
        RECT 107.590 -66.350 107.760 -66.180 ;
        RECT 108.990 -64.230 109.160 -64.060 ;
        RECT 115.580 -64.220 115.750 -64.050 ;
        RECT 108.030 -67.070 108.200 -66.900 ;
        RECT 109.040 -64.840 109.210 -64.670 ;
        RECT 115.530 -64.850 115.700 -64.680 ;
        RECT 115.580 -66.280 115.750 -66.110 ;
        RECT 109.390 -67.080 109.560 -66.910 ;
        RECT 115.180 -67.080 115.350 -66.910 ;
        RECT 115.570 -68.870 115.740 -68.700 ;
        RECT 115.970 -71.010 116.140 -70.840 ;
        RECT 116.570 -67.080 116.740 -66.910 ;
        RECT 117.010 -64.820 117.180 -64.650 ;
        RECT 117.010 -65.530 117.180 -65.360 ;
        RECT 117.970 -65.530 118.140 -65.360 ;
        RECT 118.500 -66.340 118.670 -66.170 ;
        RECT 137.330 -61.160 137.500 -60.990 ;
        RECT 139.120 -61.150 139.290 -60.980 ;
        RECT 137.790 -63.390 137.960 -63.220 ;
        RECT 140.880 -61.130 141.050 -60.960 ;
        RECT 141.990 -61.140 142.160 -60.970 ;
        RECT 119.770 -63.820 119.940 -63.650 ;
        RECT 128.570 -63.830 128.740 -63.660 ;
        RECT 119.460 -64.810 119.630 -64.640 ;
        RECT 119.460 -66.350 119.630 -66.180 ;
        RECT 120.860 -64.230 121.030 -64.060 ;
        RECT 127.450 -64.220 127.620 -64.050 ;
        RECT 119.900 -67.070 120.070 -66.900 ;
        RECT 120.910 -64.840 121.080 -64.670 ;
        RECT 127.400 -64.850 127.570 -64.680 ;
        RECT 127.450 -66.280 127.620 -66.110 ;
        RECT 121.260 -67.080 121.430 -66.910 ;
        RECT 127.050 -67.080 127.220 -66.910 ;
        RECT 127.440 -68.870 127.610 -68.700 ;
        RECT 127.840 -71.010 128.010 -70.840 ;
        RECT 128.440 -67.080 128.610 -66.910 ;
        RECT 128.880 -64.820 129.050 -64.650 ;
        RECT 128.880 -65.530 129.050 -65.360 ;
        RECT 129.840 -65.530 130.010 -65.360 ;
        RECT 130.370 -66.340 130.540 -66.170 ;
        RECT 131.640 -63.820 131.810 -63.650 ;
        RECT 137.580 -63.830 137.750 -63.660 ;
        RECT 131.330 -64.810 131.500 -64.640 ;
        RECT 131.330 -66.350 131.500 -66.180 ;
        RECT 132.730 -64.230 132.900 -64.060 ;
        RECT 136.460 -64.220 136.630 -64.050 ;
        RECT 131.770 -67.070 131.940 -66.900 ;
        RECT 132.780 -64.840 132.950 -64.670 ;
        RECT 136.410 -64.850 136.580 -64.680 ;
        RECT 136.460 -66.280 136.630 -66.110 ;
        RECT 133.130 -67.080 133.300 -66.910 ;
        RECT 136.060 -67.080 136.230 -66.910 ;
        RECT 136.450 -68.870 136.620 -68.700 ;
        RECT 136.850 -71.010 137.020 -70.840 ;
        RECT 137.450 -67.080 137.620 -66.910 ;
        RECT 137.890 -64.820 138.060 -64.650 ;
        RECT 137.890 -65.530 138.060 -65.360 ;
        RECT 138.850 -65.530 139.020 -65.360 ;
        RECT 139.380 -66.340 139.550 -66.170 ;
        RECT 140.650 -63.820 140.820 -63.650 ;
        RECT 140.340 -64.810 140.510 -64.640 ;
        RECT 140.340 -66.350 140.510 -66.180 ;
        RECT 141.740 -64.230 141.910 -64.060 ;
        RECT 140.780 -67.070 140.950 -66.900 ;
        RECT 141.790 -64.840 141.960 -64.670 ;
        RECT 142.140 -67.080 142.310 -66.910 ;
        RECT -32.870 -72.500 -32.700 -72.330 ;
        RECT -21.370 -72.500 -21.200 -72.330 ;
        RECT -9.550 -72.500 -9.380 -72.330 ;
        RECT 2.260 -72.500 2.430 -72.330 ;
        RECT 14.070 -72.500 14.240 -72.330 ;
        RECT 25.890 -72.500 26.060 -72.330 ;
        RECT 37.710 -72.500 37.880 -72.330 ;
        RECT 49.530 -72.500 49.700 -72.330 ;
        RECT 61.350 -72.500 61.520 -72.330 ;
        RECT 73.170 -72.500 73.340 -72.330 ;
        RECT 84.990 -72.500 85.160 -72.330 ;
        RECT 96.830 -72.500 97.000 -72.330 ;
        RECT 108.670 -72.500 108.840 -72.330 ;
        RECT 120.540 -72.500 120.710 -72.330 ;
        RECT 132.410 -72.500 132.580 -72.330 ;
        RECT 141.420 -72.500 141.590 -72.330 ;
        RECT -37.440 -73.900 -37.270 -73.730 ;
        RECT -37.840 -76.040 -37.670 -75.870 ;
        RECT -38.230 -77.830 -38.060 -77.660 ;
        RECT -37.880 -80.060 -37.710 -79.890 ;
        RECT -36.840 -77.830 -36.670 -77.660 ;
        RECT -37.830 -80.690 -37.660 -80.520 ;
        RECT -36.400 -79.380 -36.230 -79.210 ;
        RECT -36.400 -80.090 -36.230 -79.920 ;
        RECT -36.710 -81.080 -36.540 -80.910 ;
        RECT -35.440 -79.380 -35.270 -79.210 ;
        RECT -34.910 -78.570 -34.740 -78.400 ;
        RECT -33.950 -78.560 -33.780 -78.390 ;
        RECT -33.950 -80.100 -33.780 -79.930 ;
        RECT -32.150 -72.910 -31.980 -72.740 ;
        RECT -25.940 -73.900 -25.770 -73.730 ;
        RECT -26.340 -76.040 -26.170 -75.870 ;
        RECT -33.510 -77.840 -33.340 -77.670 ;
        RECT -32.150 -77.830 -31.980 -77.660 ;
        RECT -26.730 -77.830 -26.560 -77.660 ;
        RECT -32.500 -80.070 -32.330 -79.900 ;
        RECT -26.380 -80.060 -26.210 -79.890 ;
        RECT -25.340 -77.830 -25.170 -77.660 ;
        RECT -32.550 -80.680 -32.380 -80.510 ;
        RECT -26.330 -80.690 -26.160 -80.520 ;
        RECT -24.900 -79.380 -24.730 -79.210 ;
        RECT -24.900 -80.090 -24.730 -79.920 ;
        RECT -33.640 -81.090 -33.470 -80.920 ;
        RECT -25.210 -81.080 -25.040 -80.910 ;
        RECT -23.940 -79.380 -23.770 -79.210 ;
        RECT -23.410 -78.570 -23.240 -78.400 ;
        RECT -36.430 -81.520 -36.260 -81.350 ;
        RECT -22.450 -78.560 -22.280 -78.390 ;
        RECT -22.450 -80.100 -22.280 -79.930 ;
        RECT -20.650 -72.900 -20.480 -72.730 ;
        RECT -14.120 -73.900 -13.950 -73.730 ;
        RECT -14.520 -76.040 -14.350 -75.870 ;
        RECT -22.010 -77.840 -21.840 -77.670 ;
        RECT -20.650 -77.830 -20.480 -77.660 ;
        RECT -14.910 -77.830 -14.740 -77.660 ;
        RECT -21.000 -80.070 -20.830 -79.900 ;
        RECT -14.560 -80.060 -14.390 -79.890 ;
        RECT -13.520 -77.830 -13.350 -77.660 ;
        RECT -21.050 -80.680 -20.880 -80.510 ;
        RECT -14.510 -80.690 -14.340 -80.520 ;
        RECT -13.080 -79.380 -12.910 -79.210 ;
        RECT -13.080 -80.090 -12.910 -79.920 ;
        RECT -22.140 -81.090 -21.970 -80.920 ;
        RECT -13.390 -81.080 -13.220 -80.910 ;
        RECT -12.120 -79.380 -11.950 -79.210 ;
        RECT -11.590 -78.570 -11.420 -78.400 ;
        RECT -36.960 -83.750 -36.790 -83.580 ;
        RECT -35.170 -83.760 -35.000 -83.590 ;
        RECT -33.410 -83.780 -33.240 -83.610 ;
        RECT -25.080 -81.520 -24.910 -81.350 ;
        RECT -10.630 -78.560 -10.460 -78.390 ;
        RECT -10.630 -80.100 -10.460 -79.930 ;
        RECT -8.830 -72.900 -8.660 -72.730 ;
        RECT -2.310 -73.900 -2.140 -73.730 ;
        RECT -2.710 -76.040 -2.540 -75.870 ;
        RECT -10.190 -77.840 -10.020 -77.670 ;
        RECT -8.830 -77.830 -8.660 -77.660 ;
        RECT -3.100 -77.830 -2.930 -77.660 ;
        RECT -9.180 -80.070 -9.010 -79.900 ;
        RECT -2.750 -80.060 -2.580 -79.890 ;
        RECT -1.710 -77.830 -1.540 -77.660 ;
        RECT -9.230 -80.680 -9.060 -80.510 ;
        RECT -2.700 -80.690 -2.530 -80.520 ;
        RECT -1.270 -79.380 -1.100 -79.210 ;
        RECT -1.270 -80.090 -1.100 -79.920 ;
        RECT -10.320 -81.090 -10.150 -80.920 ;
        RECT -1.580 -81.080 -1.410 -80.910 ;
        RECT -0.310 -79.380 -0.140 -79.210 ;
        RECT 0.220 -78.570 0.390 -78.400 ;
        RECT -32.340 -83.760 -32.170 -83.590 ;
        RECT -25.460 -83.750 -25.290 -83.580 ;
        RECT -23.670 -83.760 -23.500 -83.590 ;
        RECT -21.910 -83.780 -21.740 -83.610 ;
        RECT -13.330 -81.520 -13.160 -81.350 ;
        RECT 1.180 -78.560 1.350 -78.390 ;
        RECT 1.180 -80.100 1.350 -79.930 ;
        RECT 2.980 -72.900 3.150 -72.730 ;
        RECT 9.500 -73.900 9.670 -73.730 ;
        RECT 9.100 -76.040 9.270 -75.870 ;
        RECT 1.620 -77.840 1.790 -77.670 ;
        RECT 2.980 -77.830 3.150 -77.660 ;
        RECT 8.710 -77.830 8.880 -77.660 ;
        RECT 2.630 -80.070 2.800 -79.900 ;
        RECT 9.060 -80.060 9.230 -79.890 ;
        RECT 10.100 -77.830 10.270 -77.660 ;
        RECT 2.580 -80.680 2.750 -80.510 ;
        RECT 9.110 -80.690 9.280 -80.520 ;
        RECT 10.540 -79.380 10.710 -79.210 ;
        RECT 10.540 -80.090 10.710 -79.920 ;
        RECT 1.490 -81.090 1.660 -80.920 ;
        RECT 10.230 -81.080 10.400 -80.910 ;
        RECT 11.500 -79.380 11.670 -79.210 ;
        RECT 12.030 -78.570 12.200 -78.400 ;
        RECT -20.840 -83.760 -20.670 -83.590 ;
        RECT -13.640 -83.750 -13.470 -83.580 ;
        RECT -11.850 -83.760 -11.680 -83.590 ;
        RECT -10.090 -83.780 -9.920 -83.610 ;
        RECT -1.510 -81.520 -1.340 -81.350 ;
        RECT 12.990 -78.560 13.160 -78.390 ;
        RECT 12.990 -80.100 13.160 -79.930 ;
        RECT 14.790 -72.900 14.960 -72.730 ;
        RECT 21.320 -73.900 21.490 -73.730 ;
        RECT 20.920 -76.040 21.090 -75.870 ;
        RECT 13.430 -77.840 13.600 -77.670 ;
        RECT 14.790 -77.830 14.960 -77.660 ;
        RECT 20.530 -77.830 20.700 -77.660 ;
        RECT 14.440 -80.070 14.610 -79.900 ;
        RECT 20.880 -80.060 21.050 -79.890 ;
        RECT 21.920 -77.830 22.090 -77.660 ;
        RECT 14.390 -80.680 14.560 -80.510 ;
        RECT 20.930 -80.690 21.100 -80.520 ;
        RECT 22.360 -79.380 22.530 -79.210 ;
        RECT 22.360 -80.090 22.530 -79.920 ;
        RECT 13.300 -81.090 13.470 -80.920 ;
        RECT 22.050 -81.080 22.220 -80.910 ;
        RECT 23.320 -79.380 23.490 -79.210 ;
        RECT 23.850 -78.570 24.020 -78.400 ;
        RECT -9.020 -83.760 -8.850 -83.590 ;
        RECT -1.830 -83.750 -1.660 -83.580 ;
        RECT -0.040 -83.760 0.130 -83.590 ;
        RECT 1.720 -83.780 1.890 -83.610 ;
        RECT 10.310 -81.520 10.480 -81.350 ;
        RECT 24.810 -78.560 24.980 -78.390 ;
        RECT 24.810 -80.100 24.980 -79.930 ;
        RECT 26.610 -72.900 26.780 -72.730 ;
        RECT 33.140 -73.900 33.310 -73.730 ;
        RECT 32.740 -76.040 32.910 -75.870 ;
        RECT 25.250 -77.840 25.420 -77.670 ;
        RECT 26.610 -77.830 26.780 -77.660 ;
        RECT 32.350 -77.830 32.520 -77.660 ;
        RECT 26.260 -80.070 26.430 -79.900 ;
        RECT 32.700 -80.060 32.870 -79.890 ;
        RECT 33.740 -77.830 33.910 -77.660 ;
        RECT 26.210 -80.680 26.380 -80.510 ;
        RECT 32.750 -80.690 32.920 -80.520 ;
        RECT 34.180 -79.380 34.350 -79.210 ;
        RECT 34.180 -80.090 34.350 -79.920 ;
        RECT 25.120 -81.090 25.290 -80.920 ;
        RECT 33.870 -81.080 34.040 -80.910 ;
        RECT 35.140 -79.380 35.310 -79.210 ;
        RECT 35.670 -78.570 35.840 -78.400 ;
        RECT 2.790 -83.760 2.960 -83.590 ;
        RECT 9.980 -83.750 10.150 -83.580 ;
        RECT 11.770 -83.760 11.940 -83.590 ;
        RECT 13.530 -83.780 13.700 -83.610 ;
        RECT 22.130 -81.520 22.300 -81.350 ;
        RECT 36.630 -78.560 36.800 -78.390 ;
        RECT 36.630 -80.100 36.800 -79.930 ;
        RECT 38.430 -72.900 38.600 -72.730 ;
        RECT 44.960 -73.900 45.130 -73.730 ;
        RECT 44.560 -76.040 44.730 -75.870 ;
        RECT 37.070 -77.840 37.240 -77.670 ;
        RECT 38.430 -77.830 38.600 -77.660 ;
        RECT 44.170 -77.830 44.340 -77.660 ;
        RECT 38.080 -80.070 38.250 -79.900 ;
        RECT 44.520 -80.060 44.690 -79.890 ;
        RECT 45.560 -77.830 45.730 -77.660 ;
        RECT 38.030 -80.680 38.200 -80.510 ;
        RECT 44.570 -80.690 44.740 -80.520 ;
        RECT 46.000 -79.380 46.170 -79.210 ;
        RECT 46.000 -80.090 46.170 -79.920 ;
        RECT 36.940 -81.090 37.110 -80.920 ;
        RECT 45.690 -81.080 45.860 -80.910 ;
        RECT 46.960 -79.380 47.130 -79.210 ;
        RECT 47.490 -78.570 47.660 -78.400 ;
        RECT 14.600 -83.760 14.770 -83.590 ;
        RECT 21.800 -83.750 21.970 -83.580 ;
        RECT 23.590 -83.760 23.760 -83.590 ;
        RECT 25.350 -83.780 25.520 -83.610 ;
        RECT 34.070 -81.520 34.240 -81.350 ;
        RECT 48.450 -78.560 48.620 -78.390 ;
        RECT 48.450 -80.100 48.620 -79.930 ;
        RECT 50.250 -72.900 50.420 -72.730 ;
        RECT 56.780 -73.900 56.950 -73.730 ;
        RECT 56.380 -76.040 56.550 -75.870 ;
        RECT 48.890 -77.840 49.060 -77.670 ;
        RECT 50.250 -77.830 50.420 -77.660 ;
        RECT 55.990 -77.830 56.160 -77.660 ;
        RECT 49.900 -80.070 50.070 -79.900 ;
        RECT 56.340 -80.060 56.510 -79.890 ;
        RECT 57.380 -77.830 57.550 -77.660 ;
        RECT 49.850 -80.680 50.020 -80.510 ;
        RECT 56.390 -80.690 56.560 -80.520 ;
        RECT 57.820 -79.380 57.990 -79.210 ;
        RECT 57.820 -80.090 57.990 -79.920 ;
        RECT 48.760 -81.090 48.930 -80.920 ;
        RECT 57.510 -81.080 57.680 -80.910 ;
        RECT 58.780 -79.380 58.950 -79.210 ;
        RECT 59.310 -78.570 59.480 -78.400 ;
        RECT 26.420 -83.760 26.590 -83.590 ;
        RECT 33.620 -83.750 33.790 -83.580 ;
        RECT 35.410 -83.760 35.580 -83.590 ;
        RECT 37.170 -83.780 37.340 -83.610 ;
        RECT 45.840 -81.520 46.010 -81.350 ;
        RECT 60.270 -78.560 60.440 -78.390 ;
        RECT 60.270 -80.100 60.440 -79.930 ;
        RECT 62.070 -72.900 62.240 -72.730 ;
        RECT 68.600 -73.900 68.770 -73.730 ;
        RECT 68.200 -76.040 68.370 -75.870 ;
        RECT 60.710 -77.840 60.880 -77.670 ;
        RECT 62.070 -77.830 62.240 -77.660 ;
        RECT 67.810 -77.830 67.980 -77.660 ;
        RECT 61.720 -80.070 61.890 -79.900 ;
        RECT 68.160 -80.060 68.330 -79.890 ;
        RECT 69.200 -77.830 69.370 -77.660 ;
        RECT 61.670 -80.680 61.840 -80.510 ;
        RECT 68.210 -80.690 68.380 -80.520 ;
        RECT 69.640 -79.380 69.810 -79.210 ;
        RECT 69.640 -80.090 69.810 -79.920 ;
        RECT 60.580 -81.090 60.750 -80.920 ;
        RECT 69.330 -81.080 69.500 -80.910 ;
        RECT 70.600 -79.380 70.770 -79.210 ;
        RECT 71.130 -78.570 71.300 -78.400 ;
        RECT 38.240 -83.760 38.410 -83.590 ;
        RECT 45.440 -83.750 45.610 -83.580 ;
        RECT 47.230 -83.760 47.400 -83.590 ;
        RECT 48.990 -83.780 49.160 -83.610 ;
        RECT 57.670 -81.520 57.840 -81.350 ;
        RECT 72.090 -78.560 72.260 -78.390 ;
        RECT 72.090 -80.100 72.260 -79.930 ;
        RECT 73.890 -72.900 74.060 -72.730 ;
        RECT 80.420 -73.900 80.590 -73.730 ;
        RECT 80.020 -76.040 80.190 -75.870 ;
        RECT 72.530 -77.840 72.700 -77.670 ;
        RECT 73.890 -77.830 74.060 -77.660 ;
        RECT 79.630 -77.830 79.800 -77.660 ;
        RECT 73.540 -80.070 73.710 -79.900 ;
        RECT 79.980 -80.060 80.150 -79.890 ;
        RECT 81.020 -77.830 81.190 -77.660 ;
        RECT 73.490 -80.680 73.660 -80.510 ;
        RECT 80.030 -80.690 80.200 -80.520 ;
        RECT 81.460 -79.380 81.630 -79.210 ;
        RECT 81.460 -80.090 81.630 -79.920 ;
        RECT 72.400 -81.090 72.570 -80.920 ;
        RECT 81.150 -81.080 81.320 -80.910 ;
        RECT 82.420 -79.380 82.590 -79.210 ;
        RECT 82.950 -78.570 83.120 -78.400 ;
        RECT 50.060 -83.760 50.230 -83.590 ;
        RECT 57.260 -83.750 57.430 -83.580 ;
        RECT 59.050 -83.760 59.220 -83.590 ;
        RECT 60.810 -83.780 60.980 -83.610 ;
        RECT 69.400 -81.520 69.570 -81.350 ;
        RECT 83.910 -78.560 84.080 -78.390 ;
        RECT 83.910 -80.100 84.080 -79.930 ;
        RECT 85.710 -72.900 85.880 -72.730 ;
        RECT 92.260 -73.900 92.430 -73.730 ;
        RECT 91.860 -76.040 92.030 -75.870 ;
        RECT 84.350 -77.840 84.520 -77.670 ;
        RECT 85.710 -77.830 85.880 -77.660 ;
        RECT 91.470 -77.830 91.640 -77.660 ;
        RECT 85.360 -80.070 85.530 -79.900 ;
        RECT 91.820 -80.060 91.990 -79.890 ;
        RECT 92.860 -77.830 93.030 -77.660 ;
        RECT 85.310 -80.680 85.480 -80.510 ;
        RECT 91.870 -80.690 92.040 -80.520 ;
        RECT 93.300 -79.380 93.470 -79.210 ;
        RECT 93.300 -80.090 93.470 -79.920 ;
        RECT 84.220 -81.090 84.390 -80.920 ;
        RECT 92.990 -81.080 93.160 -80.910 ;
        RECT 94.260 -79.380 94.430 -79.210 ;
        RECT 94.790 -78.570 94.960 -78.400 ;
        RECT 61.880 -83.760 62.050 -83.590 ;
        RECT 69.080 -83.750 69.250 -83.580 ;
        RECT 70.870 -83.760 71.040 -83.590 ;
        RECT 72.630 -83.780 72.800 -83.610 ;
        RECT 81.230 -81.520 81.400 -81.350 ;
        RECT 95.750 -78.560 95.920 -78.390 ;
        RECT 95.750 -80.100 95.920 -79.930 ;
        RECT 97.550 -72.900 97.720 -72.730 ;
        RECT 104.100 -73.900 104.270 -73.730 ;
        RECT 103.700 -76.040 103.870 -75.870 ;
        RECT 96.190 -77.840 96.360 -77.670 ;
        RECT 97.550 -77.830 97.720 -77.660 ;
        RECT 103.310 -77.830 103.480 -77.660 ;
        RECT 97.200 -80.070 97.370 -79.900 ;
        RECT 103.660 -80.060 103.830 -79.890 ;
        RECT 104.700 -77.830 104.870 -77.660 ;
        RECT 97.150 -80.680 97.320 -80.510 ;
        RECT 103.710 -80.690 103.880 -80.520 ;
        RECT 105.140 -79.380 105.310 -79.210 ;
        RECT 105.140 -80.090 105.310 -79.920 ;
        RECT 96.060 -81.090 96.230 -80.920 ;
        RECT 104.830 -81.080 105.000 -80.910 ;
        RECT 106.100 -79.380 106.270 -79.210 ;
        RECT 106.630 -78.570 106.800 -78.400 ;
        RECT 73.700 -83.760 73.870 -83.590 ;
        RECT 80.900 -83.750 81.070 -83.580 ;
        RECT 82.690 -83.760 82.860 -83.590 ;
        RECT 84.450 -83.780 84.620 -83.610 ;
        RECT 93.060 -81.520 93.230 -81.350 ;
        RECT 107.590 -78.560 107.760 -78.390 ;
        RECT 107.590 -80.100 107.760 -79.930 ;
        RECT 109.390 -72.900 109.560 -72.730 ;
        RECT 115.970 -73.900 116.140 -73.730 ;
        RECT 115.570 -76.040 115.740 -75.870 ;
        RECT 108.030 -77.840 108.200 -77.670 ;
        RECT 109.390 -77.830 109.560 -77.660 ;
        RECT 115.180 -77.830 115.350 -77.660 ;
        RECT 109.040 -80.070 109.210 -79.900 ;
        RECT 115.530 -80.060 115.700 -79.890 ;
        RECT 116.570 -77.830 116.740 -77.660 ;
        RECT 108.990 -80.680 109.160 -80.510 ;
        RECT 115.580 -80.690 115.750 -80.520 ;
        RECT 117.010 -79.380 117.180 -79.210 ;
        RECT 117.010 -80.090 117.180 -79.920 ;
        RECT 107.900 -81.090 108.070 -80.920 ;
        RECT 116.700 -81.080 116.870 -80.910 ;
        RECT 117.970 -79.380 118.140 -79.210 ;
        RECT 118.500 -78.570 118.670 -78.400 ;
        RECT 85.520 -83.760 85.690 -83.590 ;
        RECT 92.740 -83.750 92.910 -83.580 ;
        RECT 94.530 -83.760 94.700 -83.590 ;
        RECT 96.290 -83.780 96.460 -83.610 ;
        RECT 104.840 -81.520 105.010 -81.350 ;
        RECT 119.460 -78.560 119.630 -78.390 ;
        RECT 119.460 -80.100 119.630 -79.930 ;
        RECT 121.260 -72.900 121.430 -72.730 ;
        RECT 127.840 -73.900 128.010 -73.730 ;
        RECT 127.440 -76.040 127.610 -75.870 ;
        RECT 119.900 -77.840 120.070 -77.670 ;
        RECT 121.260 -77.830 121.430 -77.660 ;
        RECT 127.050 -77.830 127.220 -77.660 ;
        RECT 120.910 -80.070 121.080 -79.900 ;
        RECT 127.400 -80.060 127.570 -79.890 ;
        RECT 128.440 -77.830 128.610 -77.660 ;
        RECT 120.860 -80.680 121.030 -80.510 ;
        RECT 127.450 -80.690 127.620 -80.520 ;
        RECT 128.880 -79.380 129.050 -79.210 ;
        RECT 128.880 -80.090 129.050 -79.920 ;
        RECT 119.770 -81.090 119.940 -80.920 ;
        RECT 128.570 -81.080 128.740 -80.910 ;
        RECT 129.840 -79.380 130.010 -79.210 ;
        RECT 130.370 -78.570 130.540 -78.400 ;
        RECT 97.360 -83.760 97.530 -83.590 ;
        RECT 104.580 -83.750 104.750 -83.580 ;
        RECT 106.370 -83.760 106.540 -83.590 ;
        RECT 108.130 -83.780 108.300 -83.610 ;
        RECT 116.780 -81.520 116.950 -81.350 ;
        RECT 131.330 -78.560 131.500 -78.390 ;
        RECT 131.330 -80.100 131.500 -79.930 ;
        RECT 133.130 -72.900 133.300 -72.730 ;
        RECT 136.850 -73.900 137.020 -73.730 ;
        RECT 136.450 -76.040 136.620 -75.870 ;
        RECT 131.770 -77.840 131.940 -77.670 ;
        RECT 133.130 -77.830 133.300 -77.660 ;
        RECT 136.060 -77.830 136.230 -77.660 ;
        RECT 132.780 -80.070 132.950 -79.900 ;
        RECT 136.410 -80.060 136.580 -79.890 ;
        RECT 137.450 -77.830 137.620 -77.660 ;
        RECT 132.730 -80.680 132.900 -80.510 ;
        RECT 136.460 -80.690 136.630 -80.520 ;
        RECT 137.890 -79.380 138.060 -79.210 ;
        RECT 137.890 -80.090 138.060 -79.920 ;
        RECT 131.640 -81.090 131.810 -80.920 ;
        RECT 137.580 -81.080 137.750 -80.910 ;
        RECT 138.850 -79.380 139.020 -79.210 ;
        RECT 139.380 -78.570 139.550 -78.400 ;
        RECT 109.200 -83.760 109.370 -83.590 ;
        RECT 116.450 -83.750 116.620 -83.580 ;
        RECT 118.240 -83.760 118.410 -83.590 ;
        RECT 120.000 -83.780 120.170 -83.610 ;
        RECT 128.730 -81.520 128.900 -81.350 ;
        RECT 140.340 -78.560 140.510 -78.390 ;
        RECT 140.340 -80.100 140.510 -79.930 ;
        RECT 142.140 -72.900 142.310 -72.730 ;
        RECT 140.780 -77.840 140.950 -77.670 ;
        RECT 142.140 -77.830 142.310 -77.660 ;
        RECT 141.790 -80.070 141.960 -79.900 ;
        RECT 141.740 -80.680 141.910 -80.510 ;
        RECT 140.650 -81.090 140.820 -80.920 ;
        RECT 121.070 -83.760 121.240 -83.590 ;
        RECT 128.320 -83.750 128.490 -83.580 ;
        RECT 130.110 -83.760 130.280 -83.590 ;
        RECT 131.870 -83.780 132.040 -83.610 ;
        RECT 137.780 -81.520 137.950 -81.350 ;
        RECT 132.940 -83.760 133.110 -83.590 ;
        RECT 137.330 -83.750 137.500 -83.580 ;
        RECT 139.120 -83.760 139.290 -83.590 ;
        RECT 140.880 -83.780 141.050 -83.610 ;
        RECT 141.950 -83.760 142.120 -83.590 ;
        RECT -37.210 -86.120 -37.040 -85.950 ;
        RECT -33.160 -86.120 -32.990 -85.950 ;
        RECT -25.710 -86.120 -25.540 -85.950 ;
        RECT -21.660 -86.120 -21.490 -85.950 ;
        RECT -13.890 -86.120 -13.720 -85.950 ;
        RECT -9.840 -86.120 -9.670 -85.950 ;
        RECT -2.080 -86.120 -1.910 -85.950 ;
        RECT 1.970 -86.120 2.140 -85.950 ;
        RECT 9.730 -86.120 9.900 -85.950 ;
        RECT 13.780 -86.120 13.950 -85.950 ;
        RECT 21.550 -86.120 21.720 -85.950 ;
        RECT 25.600 -86.120 25.770 -85.950 ;
        RECT 33.370 -86.120 33.540 -85.950 ;
        RECT 37.420 -86.120 37.590 -85.950 ;
        RECT 45.190 -86.120 45.360 -85.950 ;
        RECT 49.240 -86.120 49.410 -85.950 ;
        RECT 57.010 -86.120 57.180 -85.950 ;
        RECT 61.060 -86.120 61.230 -85.950 ;
        RECT 68.830 -86.120 69.000 -85.950 ;
        RECT 72.880 -86.120 73.050 -85.950 ;
        RECT 80.650 -86.120 80.820 -85.950 ;
        RECT 84.700 -86.120 84.870 -85.950 ;
        RECT 92.490 -86.120 92.660 -85.950 ;
        RECT 96.540 -86.120 96.710 -85.950 ;
        RECT 104.330 -86.120 104.500 -85.950 ;
        RECT 108.380 -86.120 108.550 -85.950 ;
        RECT 116.200 -86.120 116.370 -85.950 ;
        RECT 120.250 -86.120 120.420 -85.950 ;
        RECT 128.070 -86.120 128.240 -85.950 ;
        RECT 132.120 -86.120 132.290 -85.950 ;
        RECT 137.080 -86.120 137.250 -85.950 ;
        RECT 141.130 -86.120 141.300 -85.950 ;
      LAYER met1 ;
        RECT 5.190 50.340 5.590 50.740 ;
        RECT 10.950 50.340 11.350 50.740 ;
        RECT 16.700 50.340 17.100 50.740 ;
        RECT 22.430 50.340 22.830 50.740 ;
        RECT 28.190 50.340 28.590 50.740 ;
        RECT 33.930 50.340 34.330 50.740 ;
        RECT 39.680 50.340 40.080 50.740 ;
        RECT 45.430 50.340 45.830 50.740 ;
        RECT 51.180 50.340 51.580 50.740 ;
        RECT 56.940 50.340 57.340 50.740 ;
        RECT 62.690 50.330 63.090 50.730 ;
        RECT 68.430 50.340 68.830 50.740 ;
        RECT 74.180 50.340 74.580 50.740 ;
        RECT 79.930 50.340 80.330 50.740 ;
        RECT 85.670 50.340 86.070 50.740 ;
        RECT 91.420 50.340 91.820 50.740 ;
        RECT 3.980 49.370 4.340 49.720 ;
        RECT 5.230 49.400 5.550 49.720 ;
        RECT 6.400 49.390 6.720 49.710 ;
        RECT 9.730 49.370 10.090 49.720 ;
        RECT 10.980 49.400 11.300 49.720 ;
        RECT 12.150 49.390 12.470 49.710 ;
        RECT 15.480 49.370 15.840 49.720 ;
        RECT 16.730 49.400 17.050 49.720 ;
        RECT 17.900 49.390 18.220 49.710 ;
        RECT 21.230 49.370 21.590 49.720 ;
        RECT 22.480 49.400 22.800 49.720 ;
        RECT 23.650 49.390 23.970 49.710 ;
        RECT 26.980 49.370 27.340 49.720 ;
        RECT 28.230 49.400 28.550 49.720 ;
        RECT 29.400 49.390 29.720 49.710 ;
        RECT 32.730 49.370 33.090 49.720 ;
        RECT 33.980 49.400 34.300 49.720 ;
        RECT 35.150 49.390 35.470 49.710 ;
        RECT 38.480 49.370 38.840 49.720 ;
        RECT 39.730 49.400 40.050 49.720 ;
        RECT 40.900 49.390 41.220 49.710 ;
        RECT 44.230 49.370 44.590 49.720 ;
        RECT 45.480 49.400 45.800 49.720 ;
        RECT 46.650 49.390 46.970 49.710 ;
        RECT 49.980 49.370 50.340 49.720 ;
        RECT 51.230 49.400 51.550 49.720 ;
        RECT 52.400 49.390 52.720 49.710 ;
        RECT 55.730 49.370 56.090 49.720 ;
        RECT 56.980 49.400 57.300 49.720 ;
        RECT 58.150 49.390 58.470 49.710 ;
        RECT 61.480 49.370 61.840 49.720 ;
        RECT 62.730 49.400 63.050 49.720 ;
        RECT 63.900 49.390 64.220 49.710 ;
        RECT 67.230 49.370 67.590 49.720 ;
        RECT 68.480 49.400 68.800 49.720 ;
        RECT 69.650 49.390 69.970 49.710 ;
        RECT 72.980 49.370 73.340 49.720 ;
        RECT 74.230 49.400 74.550 49.720 ;
        RECT 75.400 49.390 75.720 49.710 ;
        RECT 78.730 49.370 79.090 49.720 ;
        RECT 79.980 49.400 80.300 49.720 ;
        RECT 81.150 49.390 81.470 49.710 ;
        RECT 84.480 49.370 84.840 49.720 ;
        RECT 85.730 49.400 86.050 49.720 ;
        RECT 86.900 49.390 87.220 49.710 ;
        RECT 90.230 49.370 90.590 49.720 ;
        RECT 91.480 49.400 91.800 49.720 ;
        RECT 92.650 49.390 92.970 49.710 ;
        RECT 1.260 48.580 1.580 48.640 ;
        RECT 1.260 48.440 94.660 48.580 ;
        RECT 1.260 48.380 1.580 48.440 ;
        RECT 2.960 47.980 3.280 48.290 ;
        RECT 3.870 47.980 4.190 48.290 ;
        RECT 7.060 48.200 7.350 48.440 ;
        RECT 5.460 47.890 5.830 48.200 ;
        RECT 8.710 47.980 9.030 48.290 ;
        RECT 9.620 47.980 9.940 48.290 ;
        RECT 12.810 48.200 13.100 48.440 ;
        RECT 11.210 47.890 11.580 48.200 ;
        RECT 14.460 47.980 14.780 48.290 ;
        RECT 15.370 47.980 15.690 48.290 ;
        RECT 18.560 48.200 18.850 48.440 ;
        RECT 16.960 47.890 17.330 48.200 ;
        RECT 20.210 47.980 20.530 48.290 ;
        RECT 21.120 47.980 21.440 48.290 ;
        RECT 24.310 48.200 24.600 48.440 ;
        RECT 22.710 47.890 23.080 48.200 ;
        RECT 25.960 47.980 26.280 48.290 ;
        RECT 26.870 47.980 27.190 48.290 ;
        RECT 30.060 48.200 30.350 48.440 ;
        RECT 28.460 47.890 28.830 48.200 ;
        RECT 31.710 47.980 32.030 48.290 ;
        RECT 32.620 47.980 32.940 48.290 ;
        RECT 35.810 48.200 36.100 48.440 ;
        RECT 34.210 47.890 34.580 48.200 ;
        RECT 37.460 47.980 37.780 48.290 ;
        RECT 38.370 47.980 38.690 48.290 ;
        RECT 41.560 48.200 41.850 48.440 ;
        RECT 39.960 47.890 40.330 48.200 ;
        RECT 43.210 47.980 43.530 48.290 ;
        RECT 44.120 47.980 44.440 48.290 ;
        RECT 47.310 48.200 47.600 48.440 ;
        RECT 45.710 47.890 46.080 48.200 ;
        RECT 48.960 47.980 49.280 48.290 ;
        RECT 49.870 47.980 50.190 48.290 ;
        RECT 53.060 48.200 53.350 48.440 ;
        RECT 51.460 47.890 51.830 48.200 ;
        RECT 54.710 47.980 55.030 48.290 ;
        RECT 55.620 47.980 55.940 48.290 ;
        RECT 58.810 48.200 59.100 48.440 ;
        RECT 57.210 47.890 57.580 48.200 ;
        RECT 60.460 47.980 60.780 48.290 ;
        RECT 61.370 47.980 61.690 48.290 ;
        RECT 64.560 48.200 64.850 48.440 ;
        RECT 62.960 47.890 63.330 48.200 ;
        RECT 66.210 47.980 66.530 48.290 ;
        RECT 67.120 47.980 67.440 48.290 ;
        RECT 70.310 48.200 70.600 48.440 ;
        RECT 68.710 47.890 69.080 48.200 ;
        RECT 71.960 47.980 72.280 48.290 ;
        RECT 72.870 47.980 73.190 48.290 ;
        RECT 76.060 48.200 76.350 48.440 ;
        RECT 74.460 47.890 74.830 48.200 ;
        RECT 77.710 47.980 78.030 48.290 ;
        RECT 78.620 47.980 78.940 48.290 ;
        RECT 81.810 48.200 82.100 48.440 ;
        RECT 80.210 47.890 80.580 48.200 ;
        RECT 83.460 47.980 83.780 48.290 ;
        RECT 84.370 47.980 84.690 48.290 ;
        RECT 87.560 48.200 87.850 48.440 ;
        RECT 85.960 47.890 86.330 48.200 ;
        RECT 89.210 47.980 89.530 48.290 ;
        RECT 90.120 47.980 90.440 48.290 ;
        RECT 93.310 48.200 93.600 48.440 ;
        RECT 91.710 47.890 92.080 48.200 ;
        RECT 1.250 47.750 1.570 47.840 ;
        RECT 2.460 47.750 2.760 47.820 ;
        RECT 8.210 47.750 8.510 47.820 ;
        RECT 13.960 47.750 14.260 47.820 ;
        RECT 19.710 47.750 20.010 47.820 ;
        RECT 25.460 47.750 25.760 47.820 ;
        RECT 31.210 47.750 31.510 47.820 ;
        RECT 36.960 47.750 37.260 47.820 ;
        RECT 42.710 47.750 43.010 47.820 ;
        RECT 48.460 47.750 48.760 47.820 ;
        RECT 54.210 47.750 54.510 47.820 ;
        RECT 59.960 47.750 60.260 47.820 ;
        RECT 65.710 47.750 66.010 47.820 ;
        RECT 71.460 47.750 71.760 47.820 ;
        RECT 77.210 47.750 77.510 47.820 ;
        RECT 82.960 47.750 83.260 47.820 ;
        RECT 88.710 47.750 89.010 47.820 ;
        RECT 1.250 47.610 94.660 47.750 ;
        RECT 1.250 47.520 1.570 47.610 ;
        RECT 2.460 47.530 2.760 47.610 ;
        RECT 8.210 47.530 8.510 47.610 ;
        RECT 13.960 47.530 14.260 47.610 ;
        RECT 19.710 47.530 20.010 47.610 ;
        RECT 25.460 47.530 25.760 47.610 ;
        RECT 31.210 47.530 31.510 47.610 ;
        RECT 36.960 47.530 37.260 47.610 ;
        RECT 42.710 47.530 43.010 47.610 ;
        RECT 48.460 47.530 48.760 47.610 ;
        RECT 54.210 47.530 54.510 47.610 ;
        RECT 59.960 47.530 60.260 47.610 ;
        RECT 65.710 47.530 66.010 47.610 ;
        RECT 71.460 47.530 71.760 47.610 ;
        RECT 77.210 47.530 77.510 47.610 ;
        RECT 82.960 47.530 83.260 47.610 ;
        RECT 88.710 47.530 89.010 47.610 ;
        RECT 1.270 46.940 1.590 46.980 ;
        RECT 8.010 46.940 8.310 47.040 ;
        RECT 13.760 46.940 14.060 47.040 ;
        RECT 19.510 46.940 19.810 47.040 ;
        RECT 25.260 46.940 25.560 47.040 ;
        RECT 31.010 46.940 31.310 47.040 ;
        RECT 36.760 46.940 37.060 47.040 ;
        RECT 42.510 46.940 42.810 47.040 ;
        RECT 48.260 46.940 48.560 47.040 ;
        RECT 54.010 46.940 54.310 47.040 ;
        RECT 59.760 46.940 60.060 47.040 ;
        RECT 65.510 46.940 65.810 47.040 ;
        RECT 71.260 46.940 71.560 47.040 ;
        RECT 77.010 46.940 77.310 47.040 ;
        RECT 82.760 46.940 83.060 47.040 ;
        RECT 88.510 46.940 88.810 47.040 ;
        RECT 94.260 46.940 94.560 47.040 ;
        RECT 1.270 46.800 94.660 46.940 ;
        RECT 1.270 46.660 1.590 46.800 ;
        RECT 8.010 46.710 8.310 46.800 ;
        RECT 13.760 46.710 14.060 46.800 ;
        RECT 19.510 46.710 19.810 46.800 ;
        RECT 25.260 46.710 25.560 46.800 ;
        RECT 31.010 46.710 31.310 46.800 ;
        RECT 36.760 46.710 37.060 46.800 ;
        RECT 42.510 46.710 42.810 46.800 ;
        RECT 48.260 46.710 48.560 46.800 ;
        RECT 54.010 46.710 54.310 46.800 ;
        RECT 59.760 46.710 60.060 46.800 ;
        RECT 65.510 46.710 65.810 46.800 ;
        RECT 71.260 46.710 71.560 46.800 ;
        RECT 77.010 46.710 77.310 46.800 ;
        RECT 82.760 46.710 83.060 46.800 ;
        RECT 88.510 46.710 88.810 46.800 ;
        RECT 94.260 46.710 94.560 46.800 ;
        RECT 3.360 46.390 3.650 46.650 ;
        RECT 1.250 46.170 1.570 46.230 ;
        RECT 3.430 46.170 3.570 46.390 ;
        RECT 4.930 46.310 5.250 46.620 ;
        RECT 6.570 46.310 6.890 46.620 ;
        RECT 7.480 46.310 7.800 46.620 ;
        RECT 9.110 46.390 9.400 46.650 ;
        RECT 9.180 46.170 9.320 46.390 ;
        RECT 10.680 46.310 11.000 46.620 ;
        RECT 12.320 46.310 12.640 46.620 ;
        RECT 13.230 46.310 13.550 46.620 ;
        RECT 14.860 46.390 15.150 46.650 ;
        RECT 14.930 46.170 15.070 46.390 ;
        RECT 16.430 46.310 16.750 46.620 ;
        RECT 18.070 46.310 18.390 46.620 ;
        RECT 18.980 46.310 19.300 46.620 ;
        RECT 20.610 46.390 20.900 46.650 ;
        RECT 20.680 46.170 20.820 46.390 ;
        RECT 22.180 46.310 22.500 46.620 ;
        RECT 23.820 46.310 24.140 46.620 ;
        RECT 24.730 46.310 25.050 46.620 ;
        RECT 26.360 46.390 26.650 46.650 ;
        RECT 26.430 46.170 26.570 46.390 ;
        RECT 27.930 46.310 28.250 46.620 ;
        RECT 29.570 46.310 29.890 46.620 ;
        RECT 30.480 46.310 30.800 46.620 ;
        RECT 32.110 46.390 32.400 46.650 ;
        RECT 32.180 46.170 32.320 46.390 ;
        RECT 33.680 46.310 34.000 46.620 ;
        RECT 35.320 46.310 35.640 46.620 ;
        RECT 36.230 46.310 36.550 46.620 ;
        RECT 37.860 46.390 38.150 46.650 ;
        RECT 37.930 46.170 38.070 46.390 ;
        RECT 39.430 46.310 39.750 46.620 ;
        RECT 41.070 46.310 41.390 46.620 ;
        RECT 41.980 46.310 42.300 46.620 ;
        RECT 43.610 46.390 43.900 46.650 ;
        RECT 43.680 46.170 43.820 46.390 ;
        RECT 45.180 46.310 45.500 46.620 ;
        RECT 46.820 46.310 47.140 46.620 ;
        RECT 47.730 46.310 48.050 46.620 ;
        RECT 49.360 46.390 49.650 46.650 ;
        RECT 49.430 46.170 49.570 46.390 ;
        RECT 50.930 46.310 51.250 46.620 ;
        RECT 52.570 46.310 52.890 46.620 ;
        RECT 53.480 46.310 53.800 46.620 ;
        RECT 55.110 46.390 55.400 46.650 ;
        RECT 55.180 46.170 55.320 46.390 ;
        RECT 56.680 46.310 57.000 46.620 ;
        RECT 58.320 46.310 58.640 46.620 ;
        RECT 59.230 46.310 59.550 46.620 ;
        RECT 60.860 46.390 61.150 46.650 ;
        RECT 60.930 46.170 61.070 46.390 ;
        RECT 62.430 46.310 62.750 46.620 ;
        RECT 64.070 46.310 64.390 46.620 ;
        RECT 64.980 46.310 65.300 46.620 ;
        RECT 66.610 46.390 66.900 46.650 ;
        RECT 66.680 46.170 66.820 46.390 ;
        RECT 68.180 46.310 68.500 46.620 ;
        RECT 69.820 46.310 70.140 46.620 ;
        RECT 70.730 46.310 71.050 46.620 ;
        RECT 72.360 46.390 72.650 46.650 ;
        RECT 72.430 46.170 72.570 46.390 ;
        RECT 73.930 46.310 74.250 46.620 ;
        RECT 75.570 46.310 75.890 46.620 ;
        RECT 76.480 46.310 76.800 46.620 ;
        RECT 78.110 46.390 78.400 46.650 ;
        RECT 78.180 46.170 78.320 46.390 ;
        RECT 79.680 46.310 80.000 46.620 ;
        RECT 81.320 46.310 81.640 46.620 ;
        RECT 82.230 46.310 82.550 46.620 ;
        RECT 83.860 46.390 84.150 46.650 ;
        RECT 83.930 46.170 84.070 46.390 ;
        RECT 85.430 46.310 85.750 46.620 ;
        RECT 87.070 46.310 87.390 46.620 ;
        RECT 87.980 46.310 88.300 46.620 ;
        RECT 89.610 46.390 89.900 46.650 ;
        RECT 89.680 46.170 89.820 46.390 ;
        RECT 91.180 46.310 91.500 46.620 ;
        RECT 92.820 46.310 93.140 46.620 ;
        RECT 93.730 46.310 94.050 46.620 ;
        RECT 1.250 46.030 94.660 46.170 ;
        RECT 1.250 45.970 1.570 46.030 ;
        RECT 2.960 45.570 3.280 45.880 ;
        RECT 3.870 45.570 4.190 45.880 ;
        RECT 7.060 45.790 7.350 46.030 ;
        RECT 5.460 45.480 5.830 45.790 ;
        RECT 8.710 45.570 9.030 45.880 ;
        RECT 9.620 45.570 9.940 45.880 ;
        RECT 12.810 45.790 13.100 46.030 ;
        RECT 11.210 45.480 11.580 45.790 ;
        RECT 14.460 45.570 14.780 45.880 ;
        RECT 15.370 45.570 15.690 45.880 ;
        RECT 18.560 45.790 18.850 46.030 ;
        RECT 16.960 45.480 17.330 45.790 ;
        RECT 20.210 45.570 20.530 45.880 ;
        RECT 21.120 45.570 21.440 45.880 ;
        RECT 24.310 45.790 24.600 46.030 ;
        RECT 22.710 45.480 23.080 45.790 ;
        RECT 25.960 45.570 26.280 45.880 ;
        RECT 26.870 45.570 27.190 45.880 ;
        RECT 30.060 45.790 30.350 46.030 ;
        RECT 28.460 45.480 28.830 45.790 ;
        RECT 31.710 45.570 32.030 45.880 ;
        RECT 32.620 45.570 32.940 45.880 ;
        RECT 35.810 45.790 36.100 46.030 ;
        RECT 34.210 45.480 34.580 45.790 ;
        RECT 37.460 45.570 37.780 45.880 ;
        RECT 38.370 45.570 38.690 45.880 ;
        RECT 41.560 45.790 41.850 46.030 ;
        RECT 39.960 45.480 40.330 45.790 ;
        RECT 43.210 45.570 43.530 45.880 ;
        RECT 44.120 45.570 44.440 45.880 ;
        RECT 47.310 45.790 47.600 46.030 ;
        RECT 45.710 45.480 46.080 45.790 ;
        RECT 48.960 45.570 49.280 45.880 ;
        RECT 49.870 45.570 50.190 45.880 ;
        RECT 53.060 45.790 53.350 46.030 ;
        RECT 51.460 45.480 51.830 45.790 ;
        RECT 54.710 45.570 55.030 45.880 ;
        RECT 55.620 45.570 55.940 45.880 ;
        RECT 58.810 45.790 59.100 46.030 ;
        RECT 57.210 45.480 57.580 45.790 ;
        RECT 60.460 45.570 60.780 45.880 ;
        RECT 61.370 45.570 61.690 45.880 ;
        RECT 64.560 45.790 64.850 46.030 ;
        RECT 62.960 45.480 63.330 45.790 ;
        RECT 66.210 45.570 66.530 45.880 ;
        RECT 67.120 45.570 67.440 45.880 ;
        RECT 70.310 45.790 70.600 46.030 ;
        RECT 68.710 45.480 69.080 45.790 ;
        RECT 71.960 45.570 72.280 45.880 ;
        RECT 72.870 45.570 73.190 45.880 ;
        RECT 76.060 45.790 76.350 46.030 ;
        RECT 74.460 45.480 74.830 45.790 ;
        RECT 77.710 45.570 78.030 45.880 ;
        RECT 78.620 45.570 78.940 45.880 ;
        RECT 81.810 45.790 82.100 46.030 ;
        RECT 80.210 45.480 80.580 45.790 ;
        RECT 83.460 45.570 83.780 45.880 ;
        RECT 84.370 45.570 84.690 45.880 ;
        RECT 87.560 45.790 87.850 46.030 ;
        RECT 85.960 45.480 86.330 45.790 ;
        RECT 89.210 45.570 89.530 45.880 ;
        RECT 90.120 45.570 90.440 45.880 ;
        RECT 93.310 45.790 93.600 46.030 ;
        RECT 91.710 45.480 92.080 45.790 ;
        RECT 1.260 45.340 1.580 45.410 ;
        RECT 2.460 45.340 2.760 45.410 ;
        RECT 8.210 45.340 8.510 45.410 ;
        RECT 13.960 45.340 14.260 45.410 ;
        RECT 19.710 45.340 20.010 45.410 ;
        RECT 25.460 45.340 25.760 45.410 ;
        RECT 31.210 45.340 31.510 45.410 ;
        RECT 36.960 45.340 37.260 45.410 ;
        RECT 42.710 45.340 43.010 45.410 ;
        RECT 48.460 45.340 48.760 45.410 ;
        RECT 54.210 45.340 54.510 45.410 ;
        RECT 59.960 45.340 60.260 45.410 ;
        RECT 65.710 45.340 66.010 45.410 ;
        RECT 71.460 45.340 71.760 45.410 ;
        RECT 77.210 45.340 77.510 45.410 ;
        RECT 82.960 45.340 83.260 45.410 ;
        RECT 88.710 45.340 89.010 45.410 ;
        RECT 1.260 45.200 94.660 45.340 ;
        RECT 1.260 45.090 1.580 45.200 ;
        RECT 2.460 45.120 2.760 45.200 ;
        RECT 8.210 45.120 8.510 45.200 ;
        RECT 13.960 45.120 14.260 45.200 ;
        RECT 19.710 45.120 20.010 45.200 ;
        RECT 25.460 45.120 25.760 45.200 ;
        RECT 31.210 45.120 31.510 45.200 ;
        RECT 36.960 45.120 37.260 45.200 ;
        RECT 42.710 45.120 43.010 45.200 ;
        RECT 48.460 45.120 48.760 45.200 ;
        RECT 54.210 45.120 54.510 45.200 ;
        RECT 59.960 45.120 60.260 45.200 ;
        RECT 65.710 45.120 66.010 45.200 ;
        RECT 71.460 45.120 71.760 45.200 ;
        RECT 77.210 45.120 77.510 45.200 ;
        RECT 82.960 45.120 83.260 45.200 ;
        RECT 88.710 45.120 89.010 45.200 ;
        RECT 1.260 44.530 1.580 44.610 ;
        RECT 8.010 44.530 8.310 44.630 ;
        RECT 13.760 44.530 14.060 44.630 ;
        RECT 19.510 44.530 19.810 44.630 ;
        RECT 25.260 44.530 25.560 44.630 ;
        RECT 31.010 44.530 31.310 44.630 ;
        RECT 36.760 44.530 37.060 44.630 ;
        RECT 42.510 44.530 42.810 44.630 ;
        RECT 48.260 44.530 48.560 44.630 ;
        RECT 54.010 44.530 54.310 44.630 ;
        RECT 59.760 44.530 60.060 44.630 ;
        RECT 65.510 44.530 65.810 44.630 ;
        RECT 71.260 44.530 71.560 44.630 ;
        RECT 77.010 44.530 77.310 44.630 ;
        RECT 82.760 44.530 83.060 44.630 ;
        RECT 88.510 44.530 88.810 44.630 ;
        RECT 94.260 44.530 94.560 44.630 ;
        RECT 1.260 44.390 94.660 44.530 ;
        RECT 1.260 44.290 1.580 44.390 ;
        RECT 8.010 44.300 8.310 44.390 ;
        RECT 13.760 44.300 14.060 44.390 ;
        RECT 19.510 44.300 19.810 44.390 ;
        RECT 25.260 44.300 25.560 44.390 ;
        RECT 31.010 44.300 31.310 44.390 ;
        RECT 36.760 44.300 37.060 44.390 ;
        RECT 42.510 44.300 42.810 44.390 ;
        RECT 48.260 44.300 48.560 44.390 ;
        RECT 54.010 44.300 54.310 44.390 ;
        RECT 59.760 44.300 60.060 44.390 ;
        RECT 65.510 44.300 65.810 44.390 ;
        RECT 71.260 44.300 71.560 44.390 ;
        RECT 77.010 44.300 77.310 44.390 ;
        RECT 82.760 44.300 83.060 44.390 ;
        RECT 88.510 44.300 88.810 44.390 ;
        RECT 94.260 44.300 94.560 44.390 ;
        RECT 3.360 43.980 3.650 44.240 ;
        RECT 1.250 43.760 1.570 43.820 ;
        RECT 3.430 43.760 3.570 43.980 ;
        RECT 4.930 43.900 5.250 44.210 ;
        RECT 6.570 43.900 6.890 44.210 ;
        RECT 7.480 43.900 7.800 44.210 ;
        RECT 9.110 43.980 9.400 44.240 ;
        RECT 9.180 43.760 9.320 43.980 ;
        RECT 10.680 43.900 11.000 44.210 ;
        RECT 12.320 43.900 12.640 44.210 ;
        RECT 13.230 43.900 13.550 44.210 ;
        RECT 14.860 43.980 15.150 44.240 ;
        RECT 14.930 43.760 15.070 43.980 ;
        RECT 16.430 43.900 16.750 44.210 ;
        RECT 18.070 43.900 18.390 44.210 ;
        RECT 18.980 43.900 19.300 44.210 ;
        RECT 20.610 43.980 20.900 44.240 ;
        RECT 20.680 43.760 20.820 43.980 ;
        RECT 22.180 43.900 22.500 44.210 ;
        RECT 23.820 43.900 24.140 44.210 ;
        RECT 24.730 43.900 25.050 44.210 ;
        RECT 26.360 43.980 26.650 44.240 ;
        RECT 26.430 43.760 26.570 43.980 ;
        RECT 27.930 43.900 28.250 44.210 ;
        RECT 29.570 43.900 29.890 44.210 ;
        RECT 30.480 43.900 30.800 44.210 ;
        RECT 32.110 43.980 32.400 44.240 ;
        RECT 32.180 43.760 32.320 43.980 ;
        RECT 33.680 43.900 34.000 44.210 ;
        RECT 35.320 43.900 35.640 44.210 ;
        RECT 36.230 43.900 36.550 44.210 ;
        RECT 37.860 43.980 38.150 44.240 ;
        RECT 37.930 43.760 38.070 43.980 ;
        RECT 39.430 43.900 39.750 44.210 ;
        RECT 41.070 43.900 41.390 44.210 ;
        RECT 41.980 43.900 42.300 44.210 ;
        RECT 43.610 43.980 43.900 44.240 ;
        RECT 43.680 43.760 43.820 43.980 ;
        RECT 45.180 43.900 45.500 44.210 ;
        RECT 46.820 43.900 47.140 44.210 ;
        RECT 47.730 43.900 48.050 44.210 ;
        RECT 49.360 43.980 49.650 44.240 ;
        RECT 49.430 43.760 49.570 43.980 ;
        RECT 50.930 43.900 51.250 44.210 ;
        RECT 52.570 43.900 52.890 44.210 ;
        RECT 53.480 43.900 53.800 44.210 ;
        RECT 55.110 43.980 55.400 44.240 ;
        RECT 55.180 43.760 55.320 43.980 ;
        RECT 56.680 43.900 57.000 44.210 ;
        RECT 58.320 43.900 58.640 44.210 ;
        RECT 59.230 43.900 59.550 44.210 ;
        RECT 60.860 43.980 61.150 44.240 ;
        RECT 60.930 43.760 61.070 43.980 ;
        RECT 62.430 43.900 62.750 44.210 ;
        RECT 64.070 43.900 64.390 44.210 ;
        RECT 64.980 43.900 65.300 44.210 ;
        RECT 66.610 43.980 66.900 44.240 ;
        RECT 66.680 43.760 66.820 43.980 ;
        RECT 68.180 43.900 68.500 44.210 ;
        RECT 69.820 43.900 70.140 44.210 ;
        RECT 70.730 43.900 71.050 44.210 ;
        RECT 72.360 43.980 72.650 44.240 ;
        RECT 72.430 43.760 72.570 43.980 ;
        RECT 73.930 43.900 74.250 44.210 ;
        RECT 75.570 43.900 75.890 44.210 ;
        RECT 76.480 43.900 76.800 44.210 ;
        RECT 78.110 43.980 78.400 44.240 ;
        RECT 78.180 43.760 78.320 43.980 ;
        RECT 79.680 43.900 80.000 44.210 ;
        RECT 81.320 43.900 81.640 44.210 ;
        RECT 82.230 43.900 82.550 44.210 ;
        RECT 83.860 43.980 84.150 44.240 ;
        RECT 83.930 43.760 84.070 43.980 ;
        RECT 85.430 43.900 85.750 44.210 ;
        RECT 87.070 43.900 87.390 44.210 ;
        RECT 87.980 43.900 88.300 44.210 ;
        RECT 89.610 43.980 89.900 44.240 ;
        RECT 89.680 43.760 89.820 43.980 ;
        RECT 91.180 43.900 91.500 44.210 ;
        RECT 92.820 43.900 93.140 44.210 ;
        RECT 93.730 43.900 94.050 44.210 ;
        RECT 1.250 43.620 94.660 43.760 ;
        RECT 1.250 43.560 1.570 43.620 ;
        RECT 7.140 43.330 7.280 43.620 ;
        RECT 12.890 43.330 13.030 43.620 ;
        RECT 18.640 43.330 18.780 43.620 ;
        RECT 24.390 43.330 24.530 43.620 ;
        RECT 30.140 43.330 30.280 43.620 ;
        RECT 35.890 43.330 36.030 43.620 ;
        RECT 41.640 43.330 41.780 43.620 ;
        RECT 47.390 43.330 47.530 43.620 ;
        RECT 53.140 43.330 53.280 43.620 ;
        RECT 58.890 43.330 59.030 43.620 ;
        RECT 64.640 43.330 64.780 43.620 ;
        RECT 70.390 43.330 70.530 43.620 ;
        RECT 76.140 43.330 76.280 43.620 ;
        RECT 81.890 43.330 82.030 43.620 ;
        RECT 87.640 43.330 87.780 43.620 ;
        RECT 93.390 43.330 93.530 43.620 ;
        RECT 7.060 43.080 7.350 43.330 ;
        RECT 12.810 43.080 13.100 43.330 ;
        RECT 18.560 43.080 18.850 43.330 ;
        RECT 24.310 43.080 24.600 43.330 ;
        RECT 30.060 43.080 30.350 43.330 ;
        RECT 35.810 43.080 36.100 43.330 ;
        RECT 41.560 43.080 41.850 43.330 ;
        RECT 47.310 43.080 47.600 43.330 ;
        RECT 53.060 43.080 53.350 43.330 ;
        RECT 58.810 43.080 59.100 43.330 ;
        RECT 64.560 43.080 64.850 43.330 ;
        RECT 70.310 43.080 70.600 43.330 ;
        RECT 76.060 43.080 76.350 43.330 ;
        RECT 81.810 43.080 82.100 43.330 ;
        RECT 87.560 43.080 87.850 43.330 ;
        RECT 93.310 43.080 93.600 43.330 ;
        RECT 2.960 42.600 3.280 42.910 ;
        RECT 3.870 42.600 4.190 42.910 ;
        RECT 5.460 42.510 5.830 42.820 ;
        RECT 8.710 42.600 9.030 42.910 ;
        RECT 9.620 42.600 9.940 42.910 ;
        RECT 11.210 42.510 11.580 42.820 ;
        RECT 14.460 42.600 14.780 42.910 ;
        RECT 15.370 42.600 15.690 42.910 ;
        RECT 16.960 42.510 17.330 42.820 ;
        RECT 20.210 42.600 20.530 42.910 ;
        RECT 21.120 42.600 21.440 42.910 ;
        RECT 22.710 42.510 23.080 42.820 ;
        RECT 25.960 42.600 26.280 42.910 ;
        RECT 26.870 42.600 27.190 42.910 ;
        RECT 28.460 42.510 28.830 42.820 ;
        RECT 31.710 42.600 32.030 42.910 ;
        RECT 32.620 42.600 32.940 42.910 ;
        RECT 34.210 42.510 34.580 42.820 ;
        RECT 37.460 42.600 37.780 42.910 ;
        RECT 38.370 42.600 38.690 42.910 ;
        RECT 39.960 42.510 40.330 42.820 ;
        RECT 43.210 42.600 43.530 42.910 ;
        RECT 44.120 42.600 44.440 42.910 ;
        RECT 45.710 42.510 46.080 42.820 ;
        RECT 48.960 42.600 49.280 42.910 ;
        RECT 49.870 42.600 50.190 42.910 ;
        RECT 51.460 42.510 51.830 42.820 ;
        RECT 54.710 42.600 55.030 42.910 ;
        RECT 55.620 42.600 55.940 42.910 ;
        RECT 57.210 42.510 57.580 42.820 ;
        RECT 60.460 42.600 60.780 42.910 ;
        RECT 61.370 42.600 61.690 42.910 ;
        RECT 62.960 42.510 63.330 42.820 ;
        RECT 66.210 42.600 66.530 42.910 ;
        RECT 67.120 42.600 67.440 42.910 ;
        RECT 68.710 42.510 69.080 42.820 ;
        RECT 71.960 42.600 72.280 42.910 ;
        RECT 72.870 42.600 73.190 42.910 ;
        RECT 74.460 42.510 74.830 42.820 ;
        RECT 77.710 42.600 78.030 42.910 ;
        RECT 78.620 42.600 78.940 42.910 ;
        RECT 80.210 42.510 80.580 42.820 ;
        RECT 83.460 42.600 83.780 42.910 ;
        RECT 84.370 42.600 84.690 42.910 ;
        RECT 85.960 42.510 86.330 42.820 ;
        RECT 89.210 42.600 89.530 42.910 ;
        RECT 90.120 42.600 90.440 42.910 ;
        RECT 91.710 42.510 92.080 42.820 ;
        RECT 1.270 42.370 1.590 42.480 ;
        RECT 2.460 42.370 2.760 42.430 ;
        RECT 8.210 42.370 8.510 42.430 ;
        RECT 13.960 42.370 14.260 42.430 ;
        RECT 19.710 42.370 20.010 42.430 ;
        RECT 25.460 42.370 25.760 42.430 ;
        RECT 31.210 42.370 31.510 42.430 ;
        RECT 36.960 42.370 37.260 42.430 ;
        RECT 42.710 42.370 43.010 42.430 ;
        RECT 48.460 42.370 48.760 42.430 ;
        RECT 54.210 42.370 54.510 42.430 ;
        RECT 59.960 42.370 60.260 42.430 ;
        RECT 65.710 42.370 66.010 42.430 ;
        RECT 71.460 42.370 71.760 42.430 ;
        RECT 77.210 42.370 77.510 42.430 ;
        RECT 82.960 42.370 83.260 42.430 ;
        RECT 88.710 42.370 89.010 42.430 ;
        RECT 1.270 42.230 94.660 42.370 ;
        RECT 1.270 42.160 1.590 42.230 ;
        RECT 2.460 42.150 2.760 42.230 ;
        RECT 8.210 42.150 8.510 42.230 ;
        RECT 13.960 42.150 14.260 42.230 ;
        RECT 19.710 42.150 20.010 42.230 ;
        RECT 25.460 42.150 25.760 42.230 ;
        RECT 31.210 42.150 31.510 42.230 ;
        RECT 36.960 42.150 37.260 42.230 ;
        RECT 42.710 42.150 43.010 42.230 ;
        RECT 48.460 42.150 48.760 42.230 ;
        RECT 54.210 42.150 54.510 42.230 ;
        RECT 59.960 42.150 60.260 42.230 ;
        RECT 65.710 42.150 66.010 42.230 ;
        RECT 71.460 42.150 71.760 42.230 ;
        RECT 77.210 42.150 77.510 42.230 ;
        RECT 82.960 42.150 83.260 42.230 ;
        RECT 88.710 42.150 89.010 42.230 ;
        RECT 1.270 41.560 1.590 41.620 ;
        RECT 8.010 41.560 8.310 41.660 ;
        RECT 13.760 41.560 14.060 41.660 ;
        RECT 19.510 41.560 19.810 41.660 ;
        RECT 25.260 41.560 25.560 41.660 ;
        RECT 31.010 41.560 31.310 41.660 ;
        RECT 36.760 41.560 37.060 41.660 ;
        RECT 42.510 41.560 42.810 41.660 ;
        RECT 48.260 41.560 48.560 41.660 ;
        RECT 54.010 41.560 54.310 41.660 ;
        RECT 59.760 41.560 60.060 41.660 ;
        RECT 65.510 41.560 65.810 41.660 ;
        RECT 71.260 41.560 71.560 41.660 ;
        RECT 77.010 41.560 77.310 41.660 ;
        RECT 82.760 41.560 83.060 41.660 ;
        RECT 88.510 41.560 88.810 41.660 ;
        RECT 94.260 41.560 94.560 41.660 ;
        RECT 1.270 41.420 94.660 41.560 ;
        RECT 1.270 41.300 1.590 41.420 ;
        RECT 8.010 41.330 8.310 41.420 ;
        RECT 13.760 41.330 14.060 41.420 ;
        RECT 19.510 41.330 19.810 41.420 ;
        RECT 25.260 41.330 25.560 41.420 ;
        RECT 31.010 41.330 31.310 41.420 ;
        RECT 36.760 41.330 37.060 41.420 ;
        RECT 42.510 41.330 42.810 41.420 ;
        RECT 48.260 41.330 48.560 41.420 ;
        RECT 54.010 41.330 54.310 41.420 ;
        RECT 59.760 41.330 60.060 41.420 ;
        RECT 65.510 41.330 65.810 41.420 ;
        RECT 71.260 41.330 71.560 41.420 ;
        RECT 77.010 41.330 77.310 41.420 ;
        RECT 82.760 41.330 83.060 41.420 ;
        RECT 88.510 41.330 88.810 41.420 ;
        RECT 94.260 41.330 94.560 41.420 ;
        RECT 3.360 41.010 3.650 41.270 ;
        RECT 1.250 40.790 1.570 40.850 ;
        RECT 3.430 40.790 3.570 41.010 ;
        RECT 4.930 40.930 5.250 41.240 ;
        RECT 6.570 40.930 6.890 41.240 ;
        RECT 7.480 40.930 7.800 41.240 ;
        RECT 9.110 41.010 9.400 41.270 ;
        RECT 9.180 40.790 9.320 41.010 ;
        RECT 10.680 40.930 11.000 41.240 ;
        RECT 12.320 40.930 12.640 41.240 ;
        RECT 13.230 40.930 13.550 41.240 ;
        RECT 14.860 41.010 15.150 41.270 ;
        RECT 14.930 40.790 15.070 41.010 ;
        RECT 16.430 40.930 16.750 41.240 ;
        RECT 18.070 40.930 18.390 41.240 ;
        RECT 18.980 40.930 19.300 41.240 ;
        RECT 20.610 41.010 20.900 41.270 ;
        RECT 20.680 40.790 20.820 41.010 ;
        RECT 22.180 40.930 22.500 41.240 ;
        RECT 23.820 40.930 24.140 41.240 ;
        RECT 24.730 40.930 25.050 41.240 ;
        RECT 26.360 41.010 26.650 41.270 ;
        RECT 26.430 40.790 26.570 41.010 ;
        RECT 27.930 40.930 28.250 41.240 ;
        RECT 29.570 40.930 29.890 41.240 ;
        RECT 30.480 40.930 30.800 41.240 ;
        RECT 32.110 41.010 32.400 41.270 ;
        RECT 32.180 40.790 32.320 41.010 ;
        RECT 33.680 40.930 34.000 41.240 ;
        RECT 35.320 40.930 35.640 41.240 ;
        RECT 36.230 40.930 36.550 41.240 ;
        RECT 37.860 41.010 38.150 41.270 ;
        RECT 37.930 40.790 38.070 41.010 ;
        RECT 39.430 40.930 39.750 41.240 ;
        RECT 41.070 40.930 41.390 41.240 ;
        RECT 41.980 40.930 42.300 41.240 ;
        RECT 43.610 41.010 43.900 41.270 ;
        RECT 43.680 40.790 43.820 41.010 ;
        RECT 45.180 40.930 45.500 41.240 ;
        RECT 46.820 40.930 47.140 41.240 ;
        RECT 47.730 40.930 48.050 41.240 ;
        RECT 49.360 41.010 49.650 41.270 ;
        RECT 49.430 40.790 49.570 41.010 ;
        RECT 50.930 40.930 51.250 41.240 ;
        RECT 52.570 40.930 52.890 41.240 ;
        RECT 53.480 40.930 53.800 41.240 ;
        RECT 55.110 41.010 55.400 41.270 ;
        RECT 55.180 40.790 55.320 41.010 ;
        RECT 56.680 40.930 57.000 41.240 ;
        RECT 58.320 40.930 58.640 41.240 ;
        RECT 59.230 40.930 59.550 41.240 ;
        RECT 60.860 41.010 61.150 41.270 ;
        RECT 60.930 40.790 61.070 41.010 ;
        RECT 62.430 40.930 62.750 41.240 ;
        RECT 64.070 40.930 64.390 41.240 ;
        RECT 64.980 40.930 65.300 41.240 ;
        RECT 66.610 41.010 66.900 41.270 ;
        RECT 66.680 40.790 66.820 41.010 ;
        RECT 68.180 40.930 68.500 41.240 ;
        RECT 69.820 40.930 70.140 41.240 ;
        RECT 70.730 40.930 71.050 41.240 ;
        RECT 72.360 41.010 72.650 41.270 ;
        RECT 72.430 40.790 72.570 41.010 ;
        RECT 73.930 40.930 74.250 41.240 ;
        RECT 75.570 40.930 75.890 41.240 ;
        RECT 76.480 40.930 76.800 41.240 ;
        RECT 78.110 41.010 78.400 41.270 ;
        RECT 78.180 40.790 78.320 41.010 ;
        RECT 79.680 40.930 80.000 41.240 ;
        RECT 81.320 40.930 81.640 41.240 ;
        RECT 82.230 40.930 82.550 41.240 ;
        RECT 83.860 41.010 84.150 41.270 ;
        RECT 83.930 40.790 84.070 41.010 ;
        RECT 85.430 40.930 85.750 41.240 ;
        RECT 87.070 40.930 87.390 41.240 ;
        RECT 87.980 40.930 88.300 41.240 ;
        RECT 89.610 41.010 89.900 41.270 ;
        RECT 89.680 40.790 89.820 41.010 ;
        RECT 91.180 40.930 91.500 41.240 ;
        RECT 92.820 40.930 93.140 41.240 ;
        RECT 93.730 40.930 94.050 41.240 ;
        RECT 1.250 40.650 94.660 40.790 ;
        RECT 1.250 40.590 1.570 40.650 ;
        RECT 2.960 40.190 3.280 40.500 ;
        RECT 3.870 40.190 4.190 40.500 ;
        RECT 7.060 40.410 7.350 40.650 ;
        RECT 5.460 40.100 5.830 40.410 ;
        RECT 8.710 40.190 9.030 40.500 ;
        RECT 9.620 40.190 9.940 40.500 ;
        RECT 12.810 40.410 13.100 40.650 ;
        RECT 11.210 40.100 11.580 40.410 ;
        RECT 14.460 40.190 14.780 40.500 ;
        RECT 15.370 40.190 15.690 40.500 ;
        RECT 18.560 40.410 18.850 40.650 ;
        RECT 16.960 40.100 17.330 40.410 ;
        RECT 20.210 40.190 20.530 40.500 ;
        RECT 21.120 40.190 21.440 40.500 ;
        RECT 24.310 40.410 24.600 40.650 ;
        RECT 22.710 40.100 23.080 40.410 ;
        RECT 25.960 40.190 26.280 40.500 ;
        RECT 26.870 40.190 27.190 40.500 ;
        RECT 30.060 40.410 30.350 40.650 ;
        RECT 28.460 40.100 28.830 40.410 ;
        RECT 31.710 40.190 32.030 40.500 ;
        RECT 32.620 40.190 32.940 40.500 ;
        RECT 35.810 40.410 36.100 40.650 ;
        RECT 34.210 40.100 34.580 40.410 ;
        RECT 37.460 40.190 37.780 40.500 ;
        RECT 38.370 40.190 38.690 40.500 ;
        RECT 41.560 40.410 41.850 40.650 ;
        RECT 39.960 40.100 40.330 40.410 ;
        RECT 43.210 40.190 43.530 40.500 ;
        RECT 44.120 40.190 44.440 40.500 ;
        RECT 47.310 40.410 47.600 40.650 ;
        RECT 45.710 40.100 46.080 40.410 ;
        RECT 48.960 40.190 49.280 40.500 ;
        RECT 49.870 40.190 50.190 40.500 ;
        RECT 53.060 40.410 53.350 40.650 ;
        RECT 51.460 40.100 51.830 40.410 ;
        RECT 54.710 40.190 55.030 40.500 ;
        RECT 55.620 40.190 55.940 40.500 ;
        RECT 58.810 40.410 59.100 40.650 ;
        RECT 57.210 40.100 57.580 40.410 ;
        RECT 60.460 40.190 60.780 40.500 ;
        RECT 61.370 40.190 61.690 40.500 ;
        RECT 64.560 40.410 64.850 40.650 ;
        RECT 62.960 40.100 63.330 40.410 ;
        RECT 66.210 40.190 66.530 40.500 ;
        RECT 67.120 40.190 67.440 40.500 ;
        RECT 70.310 40.410 70.600 40.650 ;
        RECT 68.710 40.100 69.080 40.410 ;
        RECT 71.960 40.190 72.280 40.500 ;
        RECT 72.870 40.190 73.190 40.500 ;
        RECT 76.060 40.410 76.350 40.650 ;
        RECT 74.460 40.100 74.830 40.410 ;
        RECT 77.710 40.190 78.030 40.500 ;
        RECT 78.620 40.190 78.940 40.500 ;
        RECT 81.810 40.410 82.100 40.650 ;
        RECT 80.210 40.100 80.580 40.410 ;
        RECT 83.460 40.190 83.780 40.500 ;
        RECT 84.370 40.190 84.690 40.500 ;
        RECT 87.560 40.410 87.850 40.650 ;
        RECT 85.960 40.100 86.330 40.410 ;
        RECT 89.210 40.190 89.530 40.500 ;
        RECT 90.120 40.190 90.440 40.500 ;
        RECT 93.310 40.410 93.600 40.650 ;
        RECT 91.710 40.100 92.080 40.410 ;
        RECT 1.270 39.960 1.590 40.050 ;
        RECT 2.460 39.960 2.760 40.030 ;
        RECT 8.210 39.960 8.510 40.030 ;
        RECT 13.960 39.960 14.260 40.030 ;
        RECT 19.710 39.960 20.010 40.030 ;
        RECT 25.460 39.960 25.760 40.030 ;
        RECT 31.210 39.960 31.510 40.030 ;
        RECT 36.960 39.960 37.260 40.030 ;
        RECT 42.710 39.960 43.010 40.030 ;
        RECT 48.460 39.960 48.760 40.030 ;
        RECT 54.210 39.960 54.510 40.030 ;
        RECT 59.960 39.960 60.260 40.030 ;
        RECT 65.710 39.960 66.010 40.030 ;
        RECT 71.460 39.960 71.760 40.030 ;
        RECT 77.210 39.960 77.510 40.030 ;
        RECT 82.960 39.960 83.260 40.030 ;
        RECT 88.710 39.960 89.010 40.030 ;
        RECT 1.270 39.820 94.660 39.960 ;
        RECT 1.270 39.730 1.590 39.820 ;
        RECT 2.460 39.740 2.760 39.820 ;
        RECT 8.210 39.740 8.510 39.820 ;
        RECT 13.960 39.740 14.260 39.820 ;
        RECT 19.710 39.740 20.010 39.820 ;
        RECT 25.460 39.740 25.760 39.820 ;
        RECT 31.210 39.740 31.510 39.820 ;
        RECT 36.960 39.740 37.260 39.820 ;
        RECT 42.710 39.740 43.010 39.820 ;
        RECT 48.460 39.740 48.760 39.820 ;
        RECT 54.210 39.740 54.510 39.820 ;
        RECT 59.960 39.740 60.260 39.820 ;
        RECT 65.710 39.740 66.010 39.820 ;
        RECT 71.460 39.740 71.760 39.820 ;
        RECT 77.210 39.740 77.510 39.820 ;
        RECT 82.960 39.740 83.260 39.820 ;
        RECT 88.710 39.740 89.010 39.820 ;
        RECT 1.270 39.150 1.590 39.210 ;
        RECT 8.010 39.150 8.310 39.250 ;
        RECT 13.760 39.150 14.060 39.250 ;
        RECT 19.510 39.150 19.810 39.250 ;
        RECT 25.260 39.150 25.560 39.250 ;
        RECT 31.010 39.150 31.310 39.250 ;
        RECT 36.760 39.150 37.060 39.250 ;
        RECT 42.510 39.150 42.810 39.250 ;
        RECT 48.260 39.150 48.560 39.250 ;
        RECT 54.010 39.150 54.310 39.250 ;
        RECT 59.760 39.150 60.060 39.250 ;
        RECT 65.510 39.150 65.810 39.250 ;
        RECT 71.260 39.150 71.560 39.250 ;
        RECT 77.010 39.150 77.310 39.250 ;
        RECT 82.760 39.150 83.060 39.250 ;
        RECT 88.510 39.150 88.810 39.250 ;
        RECT 94.260 39.150 94.560 39.250 ;
        RECT 1.270 39.010 94.660 39.150 ;
        RECT 1.270 38.890 1.590 39.010 ;
        RECT 8.010 38.920 8.310 39.010 ;
        RECT 13.760 38.920 14.060 39.010 ;
        RECT 19.510 38.920 19.810 39.010 ;
        RECT 25.260 38.920 25.560 39.010 ;
        RECT 31.010 38.920 31.310 39.010 ;
        RECT 36.760 38.920 37.060 39.010 ;
        RECT 42.510 38.920 42.810 39.010 ;
        RECT 48.260 38.920 48.560 39.010 ;
        RECT 54.010 38.920 54.310 39.010 ;
        RECT 59.760 38.920 60.060 39.010 ;
        RECT 65.510 38.920 65.810 39.010 ;
        RECT 71.260 38.920 71.560 39.010 ;
        RECT 77.010 38.920 77.310 39.010 ;
        RECT 82.760 38.920 83.060 39.010 ;
        RECT 88.510 38.920 88.810 39.010 ;
        RECT 94.260 38.920 94.560 39.010 ;
        RECT 3.360 38.600 3.650 38.860 ;
        RECT 1.260 38.380 1.580 38.440 ;
        RECT 3.430 38.380 3.570 38.600 ;
        RECT 4.930 38.520 5.250 38.830 ;
        RECT 6.570 38.520 6.890 38.830 ;
        RECT 7.480 38.520 7.800 38.830 ;
        RECT 9.110 38.600 9.400 38.860 ;
        RECT 9.180 38.380 9.320 38.600 ;
        RECT 10.680 38.520 11.000 38.830 ;
        RECT 12.320 38.520 12.640 38.830 ;
        RECT 13.230 38.520 13.550 38.830 ;
        RECT 14.860 38.600 15.150 38.860 ;
        RECT 14.930 38.380 15.070 38.600 ;
        RECT 16.430 38.520 16.750 38.830 ;
        RECT 18.070 38.520 18.390 38.830 ;
        RECT 18.980 38.520 19.300 38.830 ;
        RECT 20.610 38.600 20.900 38.860 ;
        RECT 20.680 38.380 20.820 38.600 ;
        RECT 22.180 38.520 22.500 38.830 ;
        RECT 23.820 38.520 24.140 38.830 ;
        RECT 24.730 38.520 25.050 38.830 ;
        RECT 26.360 38.600 26.650 38.860 ;
        RECT 26.430 38.380 26.570 38.600 ;
        RECT 27.930 38.520 28.250 38.830 ;
        RECT 29.570 38.520 29.890 38.830 ;
        RECT 30.480 38.520 30.800 38.830 ;
        RECT 32.110 38.600 32.400 38.860 ;
        RECT 32.180 38.380 32.320 38.600 ;
        RECT 33.680 38.520 34.000 38.830 ;
        RECT 35.320 38.520 35.640 38.830 ;
        RECT 36.230 38.520 36.550 38.830 ;
        RECT 37.860 38.600 38.150 38.860 ;
        RECT 37.930 38.380 38.070 38.600 ;
        RECT 39.430 38.520 39.750 38.830 ;
        RECT 41.070 38.520 41.390 38.830 ;
        RECT 41.980 38.520 42.300 38.830 ;
        RECT 43.610 38.600 43.900 38.860 ;
        RECT 43.680 38.380 43.820 38.600 ;
        RECT 45.180 38.520 45.500 38.830 ;
        RECT 46.820 38.520 47.140 38.830 ;
        RECT 47.730 38.520 48.050 38.830 ;
        RECT 49.360 38.600 49.650 38.860 ;
        RECT 49.430 38.380 49.570 38.600 ;
        RECT 50.930 38.520 51.250 38.830 ;
        RECT 52.570 38.520 52.890 38.830 ;
        RECT 53.480 38.520 53.800 38.830 ;
        RECT 55.110 38.600 55.400 38.860 ;
        RECT 55.180 38.380 55.320 38.600 ;
        RECT 56.680 38.520 57.000 38.830 ;
        RECT 58.320 38.520 58.640 38.830 ;
        RECT 59.230 38.520 59.550 38.830 ;
        RECT 60.860 38.600 61.150 38.860 ;
        RECT 60.930 38.380 61.070 38.600 ;
        RECT 62.430 38.520 62.750 38.830 ;
        RECT 64.070 38.520 64.390 38.830 ;
        RECT 64.980 38.520 65.300 38.830 ;
        RECT 66.610 38.600 66.900 38.860 ;
        RECT 66.680 38.380 66.820 38.600 ;
        RECT 68.180 38.520 68.500 38.830 ;
        RECT 69.820 38.520 70.140 38.830 ;
        RECT 70.730 38.520 71.050 38.830 ;
        RECT 72.360 38.600 72.650 38.860 ;
        RECT 72.430 38.380 72.570 38.600 ;
        RECT 73.930 38.520 74.250 38.830 ;
        RECT 75.570 38.520 75.890 38.830 ;
        RECT 76.480 38.520 76.800 38.830 ;
        RECT 78.110 38.600 78.400 38.860 ;
        RECT 78.180 38.380 78.320 38.600 ;
        RECT 79.680 38.520 80.000 38.830 ;
        RECT 81.320 38.520 81.640 38.830 ;
        RECT 82.230 38.520 82.550 38.830 ;
        RECT 83.860 38.600 84.150 38.860 ;
        RECT 83.930 38.380 84.070 38.600 ;
        RECT 85.430 38.520 85.750 38.830 ;
        RECT 87.070 38.520 87.390 38.830 ;
        RECT 87.980 38.520 88.300 38.830 ;
        RECT 89.610 38.600 89.900 38.860 ;
        RECT 89.680 38.380 89.820 38.600 ;
        RECT 91.180 38.520 91.500 38.830 ;
        RECT 92.820 38.520 93.140 38.830 ;
        RECT 93.730 38.520 94.050 38.830 ;
        RECT 1.260 38.240 94.660 38.380 ;
        RECT 1.260 38.180 1.580 38.240 ;
        RECT 2.960 37.780 3.280 38.090 ;
        RECT 3.870 37.780 4.190 38.090 ;
        RECT 7.060 38.000 7.350 38.240 ;
        RECT 5.460 37.690 5.830 38.000 ;
        RECT 8.710 37.780 9.030 38.090 ;
        RECT 9.620 37.780 9.940 38.090 ;
        RECT 12.810 38.000 13.100 38.240 ;
        RECT 11.210 37.690 11.580 38.000 ;
        RECT 14.460 37.780 14.780 38.090 ;
        RECT 15.370 37.780 15.690 38.090 ;
        RECT 18.560 38.000 18.850 38.240 ;
        RECT 16.960 37.690 17.330 38.000 ;
        RECT 20.210 37.780 20.530 38.090 ;
        RECT 21.120 37.780 21.440 38.090 ;
        RECT 24.310 38.000 24.600 38.240 ;
        RECT 22.710 37.690 23.080 38.000 ;
        RECT 25.960 37.780 26.280 38.090 ;
        RECT 26.870 37.780 27.190 38.090 ;
        RECT 30.060 38.000 30.350 38.240 ;
        RECT 28.460 37.690 28.830 38.000 ;
        RECT 31.710 37.780 32.030 38.090 ;
        RECT 32.620 37.780 32.940 38.090 ;
        RECT 35.810 38.000 36.100 38.240 ;
        RECT 34.210 37.690 34.580 38.000 ;
        RECT 37.460 37.780 37.780 38.090 ;
        RECT 38.370 37.780 38.690 38.090 ;
        RECT 41.560 38.000 41.850 38.240 ;
        RECT 39.960 37.690 40.330 38.000 ;
        RECT 43.210 37.780 43.530 38.090 ;
        RECT 44.120 37.780 44.440 38.090 ;
        RECT 47.310 38.000 47.600 38.240 ;
        RECT 45.710 37.690 46.080 38.000 ;
        RECT 48.960 37.780 49.280 38.090 ;
        RECT 49.870 37.780 50.190 38.090 ;
        RECT 53.060 38.000 53.350 38.240 ;
        RECT 51.460 37.690 51.830 38.000 ;
        RECT 54.710 37.780 55.030 38.090 ;
        RECT 55.620 37.780 55.940 38.090 ;
        RECT 58.810 38.000 59.100 38.240 ;
        RECT 57.210 37.690 57.580 38.000 ;
        RECT 60.460 37.780 60.780 38.090 ;
        RECT 61.370 37.780 61.690 38.090 ;
        RECT 64.560 38.000 64.850 38.240 ;
        RECT 62.960 37.690 63.330 38.000 ;
        RECT 66.210 37.780 66.530 38.090 ;
        RECT 67.120 37.780 67.440 38.090 ;
        RECT 70.310 38.000 70.600 38.240 ;
        RECT 68.710 37.690 69.080 38.000 ;
        RECT 71.960 37.780 72.280 38.090 ;
        RECT 72.870 37.780 73.190 38.090 ;
        RECT 76.060 38.000 76.350 38.240 ;
        RECT 74.460 37.690 74.830 38.000 ;
        RECT 77.710 37.780 78.030 38.090 ;
        RECT 78.620 37.780 78.940 38.090 ;
        RECT 81.810 38.000 82.100 38.240 ;
        RECT 80.210 37.690 80.580 38.000 ;
        RECT 83.460 37.780 83.780 38.090 ;
        RECT 84.370 37.780 84.690 38.090 ;
        RECT 87.560 38.000 87.850 38.240 ;
        RECT 85.960 37.690 86.330 38.000 ;
        RECT 89.210 37.780 89.530 38.090 ;
        RECT 90.120 37.780 90.440 38.090 ;
        RECT 93.310 38.000 93.600 38.240 ;
        RECT 91.710 37.690 92.080 38.000 ;
        RECT 3.360 36.190 3.650 36.450 ;
        RECT 1.260 35.970 1.580 36.030 ;
        RECT 3.430 35.970 3.570 36.190 ;
        RECT 4.930 36.110 5.250 36.420 ;
        RECT 6.570 36.110 6.890 36.420 ;
        RECT 7.480 36.110 7.800 36.420 ;
        RECT 9.110 36.190 9.400 36.450 ;
        RECT 9.180 35.970 9.320 36.190 ;
        RECT 10.680 36.110 11.000 36.420 ;
        RECT 12.320 36.110 12.640 36.420 ;
        RECT 13.230 36.110 13.550 36.420 ;
        RECT 14.860 36.190 15.150 36.450 ;
        RECT 14.930 35.970 15.070 36.190 ;
        RECT 16.430 36.110 16.750 36.420 ;
        RECT 18.070 36.110 18.390 36.420 ;
        RECT 18.980 36.110 19.300 36.420 ;
        RECT 20.610 36.190 20.900 36.450 ;
        RECT 20.680 35.970 20.820 36.190 ;
        RECT 22.180 36.110 22.500 36.420 ;
        RECT 23.820 36.110 24.140 36.420 ;
        RECT 24.730 36.110 25.050 36.420 ;
        RECT 26.360 36.190 26.650 36.450 ;
        RECT 26.430 35.970 26.570 36.190 ;
        RECT 27.930 36.110 28.250 36.420 ;
        RECT 29.570 36.110 29.890 36.420 ;
        RECT 30.480 36.110 30.800 36.420 ;
        RECT 32.110 36.190 32.400 36.450 ;
        RECT 32.180 35.970 32.320 36.190 ;
        RECT 33.680 36.110 34.000 36.420 ;
        RECT 35.320 36.110 35.640 36.420 ;
        RECT 36.230 36.110 36.550 36.420 ;
        RECT 37.860 36.190 38.150 36.450 ;
        RECT 37.930 35.970 38.070 36.190 ;
        RECT 39.430 36.110 39.750 36.420 ;
        RECT 41.070 36.110 41.390 36.420 ;
        RECT 41.980 36.110 42.300 36.420 ;
        RECT 43.610 36.190 43.900 36.450 ;
        RECT 43.680 35.970 43.820 36.190 ;
        RECT 45.180 36.110 45.500 36.420 ;
        RECT 46.820 36.110 47.140 36.420 ;
        RECT 47.730 36.110 48.050 36.420 ;
        RECT 49.360 36.190 49.650 36.450 ;
        RECT 49.430 35.970 49.570 36.190 ;
        RECT 50.930 36.110 51.250 36.420 ;
        RECT 52.570 36.110 52.890 36.420 ;
        RECT 53.480 36.110 53.800 36.420 ;
        RECT 55.110 36.190 55.400 36.450 ;
        RECT 55.180 35.970 55.320 36.190 ;
        RECT 56.680 36.110 57.000 36.420 ;
        RECT 58.320 36.110 58.640 36.420 ;
        RECT 59.230 36.110 59.550 36.420 ;
        RECT 60.860 36.190 61.150 36.450 ;
        RECT 60.930 35.970 61.070 36.190 ;
        RECT 62.430 36.110 62.750 36.420 ;
        RECT 64.070 36.110 64.390 36.420 ;
        RECT 64.980 36.110 65.300 36.420 ;
        RECT 66.610 36.190 66.900 36.450 ;
        RECT 66.680 35.970 66.820 36.190 ;
        RECT 68.180 36.110 68.500 36.420 ;
        RECT 69.820 36.110 70.140 36.420 ;
        RECT 70.730 36.110 71.050 36.420 ;
        RECT 72.360 36.190 72.650 36.450 ;
        RECT 72.430 35.970 72.570 36.190 ;
        RECT 73.930 36.110 74.250 36.420 ;
        RECT 75.570 36.110 75.890 36.420 ;
        RECT 76.480 36.110 76.800 36.420 ;
        RECT 78.110 36.190 78.400 36.450 ;
        RECT 78.180 35.970 78.320 36.190 ;
        RECT 79.680 36.110 80.000 36.420 ;
        RECT 81.320 36.110 81.640 36.420 ;
        RECT 82.230 36.110 82.550 36.420 ;
        RECT 83.860 36.190 84.150 36.450 ;
        RECT 83.930 35.970 84.070 36.190 ;
        RECT 85.430 36.110 85.750 36.420 ;
        RECT 87.070 36.110 87.390 36.420 ;
        RECT 87.980 36.110 88.300 36.420 ;
        RECT 89.610 36.190 89.900 36.450 ;
        RECT 89.680 35.970 89.820 36.190 ;
        RECT 91.180 36.110 91.500 36.420 ;
        RECT 92.820 36.110 93.140 36.420 ;
        RECT 93.730 36.110 94.050 36.420 ;
        RECT 1.260 35.830 94.660 35.970 ;
        RECT 1.260 35.770 1.580 35.830 ;
        RECT 2.960 35.370 3.280 35.680 ;
        RECT 3.870 35.370 4.190 35.680 ;
        RECT 7.060 35.590 7.350 35.830 ;
        RECT 5.460 35.280 5.830 35.590 ;
        RECT 8.710 35.370 9.030 35.680 ;
        RECT 9.620 35.370 9.940 35.680 ;
        RECT 12.810 35.590 13.100 35.830 ;
        RECT 11.210 35.280 11.580 35.590 ;
        RECT 14.460 35.370 14.780 35.680 ;
        RECT 15.370 35.370 15.690 35.680 ;
        RECT 18.560 35.590 18.850 35.830 ;
        RECT 16.960 35.280 17.330 35.590 ;
        RECT 20.210 35.370 20.530 35.680 ;
        RECT 21.120 35.370 21.440 35.680 ;
        RECT 24.310 35.590 24.600 35.830 ;
        RECT 22.710 35.280 23.080 35.590 ;
        RECT 25.960 35.370 26.280 35.680 ;
        RECT 26.870 35.370 27.190 35.680 ;
        RECT 30.060 35.590 30.350 35.830 ;
        RECT 28.460 35.280 28.830 35.590 ;
        RECT 31.710 35.370 32.030 35.680 ;
        RECT 32.620 35.370 32.940 35.680 ;
        RECT 35.810 35.590 36.100 35.830 ;
        RECT 34.210 35.280 34.580 35.590 ;
        RECT 37.460 35.370 37.780 35.680 ;
        RECT 38.370 35.370 38.690 35.680 ;
        RECT 41.560 35.590 41.850 35.830 ;
        RECT 39.960 35.280 40.330 35.590 ;
        RECT 43.210 35.370 43.530 35.680 ;
        RECT 44.120 35.370 44.440 35.680 ;
        RECT 47.310 35.590 47.600 35.830 ;
        RECT 45.710 35.280 46.080 35.590 ;
        RECT 48.960 35.370 49.280 35.680 ;
        RECT 49.870 35.370 50.190 35.680 ;
        RECT 53.060 35.590 53.350 35.830 ;
        RECT 51.460 35.280 51.830 35.590 ;
        RECT 54.710 35.370 55.030 35.680 ;
        RECT 55.620 35.370 55.940 35.680 ;
        RECT 58.810 35.590 59.100 35.830 ;
        RECT 57.210 35.280 57.580 35.590 ;
        RECT 60.460 35.370 60.780 35.680 ;
        RECT 61.370 35.370 61.690 35.680 ;
        RECT 64.560 35.590 64.850 35.830 ;
        RECT 62.960 35.280 63.330 35.590 ;
        RECT 66.210 35.370 66.530 35.680 ;
        RECT 67.120 35.370 67.440 35.680 ;
        RECT 70.310 35.590 70.600 35.830 ;
        RECT 68.710 35.280 69.080 35.590 ;
        RECT 71.960 35.370 72.280 35.680 ;
        RECT 72.870 35.370 73.190 35.680 ;
        RECT 76.060 35.590 76.350 35.830 ;
        RECT 74.460 35.280 74.830 35.590 ;
        RECT 77.710 35.370 78.030 35.680 ;
        RECT 78.620 35.370 78.940 35.680 ;
        RECT 81.810 35.590 82.100 35.830 ;
        RECT 80.210 35.280 80.580 35.590 ;
        RECT 83.460 35.370 83.780 35.680 ;
        RECT 84.370 35.370 84.690 35.680 ;
        RECT 87.560 35.590 87.850 35.830 ;
        RECT 85.960 35.280 86.330 35.590 ;
        RECT 89.210 35.370 89.530 35.680 ;
        RECT 90.120 35.370 90.440 35.680 ;
        RECT 93.310 35.590 93.600 35.830 ;
        RECT 91.710 35.280 92.080 35.590 ;
        RECT 3.360 33.780 3.650 34.040 ;
        RECT 1.260 33.560 1.580 33.620 ;
        RECT 3.430 33.560 3.570 33.780 ;
        RECT 4.930 33.700 5.250 34.010 ;
        RECT 6.570 33.700 6.890 34.010 ;
        RECT 7.480 33.700 7.800 34.010 ;
        RECT 9.110 33.780 9.400 34.040 ;
        RECT 9.180 33.560 9.320 33.780 ;
        RECT 10.680 33.700 11.000 34.010 ;
        RECT 12.320 33.700 12.640 34.010 ;
        RECT 13.230 33.700 13.550 34.010 ;
        RECT 14.860 33.780 15.150 34.040 ;
        RECT 14.930 33.560 15.070 33.780 ;
        RECT 16.430 33.700 16.750 34.010 ;
        RECT 18.070 33.700 18.390 34.010 ;
        RECT 18.980 33.700 19.300 34.010 ;
        RECT 20.610 33.780 20.900 34.040 ;
        RECT 20.680 33.560 20.820 33.780 ;
        RECT 22.180 33.700 22.500 34.010 ;
        RECT 23.820 33.700 24.140 34.010 ;
        RECT 24.730 33.700 25.050 34.010 ;
        RECT 26.360 33.780 26.650 34.040 ;
        RECT 26.430 33.560 26.570 33.780 ;
        RECT 27.930 33.700 28.250 34.010 ;
        RECT 29.570 33.700 29.890 34.010 ;
        RECT 30.480 33.700 30.800 34.010 ;
        RECT 32.110 33.780 32.400 34.040 ;
        RECT 32.180 33.560 32.320 33.780 ;
        RECT 33.680 33.700 34.000 34.010 ;
        RECT 35.320 33.700 35.640 34.010 ;
        RECT 36.230 33.700 36.550 34.010 ;
        RECT 37.860 33.780 38.150 34.040 ;
        RECT 37.930 33.560 38.070 33.780 ;
        RECT 39.430 33.700 39.750 34.010 ;
        RECT 41.070 33.700 41.390 34.010 ;
        RECT 41.980 33.700 42.300 34.010 ;
        RECT 43.610 33.780 43.900 34.040 ;
        RECT 43.680 33.560 43.820 33.780 ;
        RECT 45.180 33.700 45.500 34.010 ;
        RECT 46.820 33.700 47.140 34.010 ;
        RECT 47.730 33.700 48.050 34.010 ;
        RECT 49.360 33.780 49.650 34.040 ;
        RECT 49.430 33.560 49.570 33.780 ;
        RECT 50.930 33.700 51.250 34.010 ;
        RECT 52.570 33.700 52.890 34.010 ;
        RECT 53.480 33.700 53.800 34.010 ;
        RECT 55.110 33.780 55.400 34.040 ;
        RECT 55.180 33.560 55.320 33.780 ;
        RECT 56.680 33.700 57.000 34.010 ;
        RECT 58.320 33.700 58.640 34.010 ;
        RECT 59.230 33.700 59.550 34.010 ;
        RECT 60.860 33.780 61.150 34.040 ;
        RECT 60.930 33.560 61.070 33.780 ;
        RECT 62.430 33.700 62.750 34.010 ;
        RECT 64.070 33.700 64.390 34.010 ;
        RECT 64.980 33.700 65.300 34.010 ;
        RECT 66.610 33.780 66.900 34.040 ;
        RECT 66.680 33.560 66.820 33.780 ;
        RECT 68.180 33.700 68.500 34.010 ;
        RECT 69.820 33.700 70.140 34.010 ;
        RECT 70.730 33.700 71.050 34.010 ;
        RECT 72.360 33.780 72.650 34.040 ;
        RECT 72.430 33.560 72.570 33.780 ;
        RECT 73.930 33.700 74.250 34.010 ;
        RECT 75.570 33.700 75.890 34.010 ;
        RECT 76.480 33.700 76.800 34.010 ;
        RECT 78.110 33.780 78.400 34.040 ;
        RECT 78.180 33.560 78.320 33.780 ;
        RECT 79.680 33.700 80.000 34.010 ;
        RECT 81.320 33.700 81.640 34.010 ;
        RECT 82.230 33.700 82.550 34.010 ;
        RECT 83.860 33.780 84.150 34.040 ;
        RECT 83.930 33.560 84.070 33.780 ;
        RECT 85.430 33.700 85.750 34.010 ;
        RECT 87.070 33.700 87.390 34.010 ;
        RECT 87.980 33.700 88.300 34.010 ;
        RECT 89.610 33.780 89.900 34.040 ;
        RECT 89.680 33.560 89.820 33.780 ;
        RECT 91.180 33.700 91.500 34.010 ;
        RECT 92.820 33.700 93.140 34.010 ;
        RECT 93.730 33.700 94.050 34.010 ;
        RECT 1.260 33.420 94.660 33.560 ;
        RECT 1.260 33.360 1.580 33.420 ;
        RECT 2.960 32.960 3.280 33.270 ;
        RECT 3.870 32.960 4.190 33.270 ;
        RECT 7.060 33.180 7.350 33.420 ;
        RECT 5.460 32.870 5.830 33.180 ;
        RECT 8.710 32.960 9.030 33.270 ;
        RECT 9.620 32.960 9.940 33.270 ;
        RECT 12.810 33.180 13.100 33.420 ;
        RECT 11.210 32.870 11.580 33.180 ;
        RECT 14.460 32.960 14.780 33.270 ;
        RECT 15.370 32.960 15.690 33.270 ;
        RECT 18.560 33.180 18.850 33.420 ;
        RECT 16.960 32.870 17.330 33.180 ;
        RECT 20.210 32.960 20.530 33.270 ;
        RECT 21.120 32.960 21.440 33.270 ;
        RECT 24.310 33.180 24.600 33.420 ;
        RECT 22.710 32.870 23.080 33.180 ;
        RECT 25.960 32.960 26.280 33.270 ;
        RECT 26.870 32.960 27.190 33.270 ;
        RECT 30.060 33.180 30.350 33.420 ;
        RECT 28.460 32.870 28.830 33.180 ;
        RECT 31.710 32.960 32.030 33.270 ;
        RECT 32.620 32.960 32.940 33.270 ;
        RECT 35.810 33.180 36.100 33.420 ;
        RECT 34.210 32.870 34.580 33.180 ;
        RECT 37.460 32.960 37.780 33.270 ;
        RECT 38.370 32.960 38.690 33.270 ;
        RECT 41.560 33.180 41.850 33.420 ;
        RECT 39.960 32.870 40.330 33.180 ;
        RECT 43.210 32.960 43.530 33.270 ;
        RECT 44.120 32.960 44.440 33.270 ;
        RECT 47.310 33.180 47.600 33.420 ;
        RECT 45.710 32.870 46.080 33.180 ;
        RECT 48.960 32.960 49.280 33.270 ;
        RECT 49.870 32.960 50.190 33.270 ;
        RECT 53.060 33.180 53.350 33.420 ;
        RECT 51.460 32.870 51.830 33.180 ;
        RECT 54.710 32.960 55.030 33.270 ;
        RECT 55.620 32.960 55.940 33.270 ;
        RECT 58.810 33.180 59.100 33.420 ;
        RECT 57.210 32.870 57.580 33.180 ;
        RECT 60.460 32.960 60.780 33.270 ;
        RECT 61.370 32.960 61.690 33.270 ;
        RECT 64.560 33.180 64.850 33.420 ;
        RECT 62.960 32.870 63.330 33.180 ;
        RECT 66.210 32.960 66.530 33.270 ;
        RECT 67.120 32.960 67.440 33.270 ;
        RECT 70.310 33.180 70.600 33.420 ;
        RECT 68.710 32.870 69.080 33.180 ;
        RECT 71.960 32.960 72.280 33.270 ;
        RECT 72.870 32.960 73.190 33.270 ;
        RECT 76.060 33.180 76.350 33.420 ;
        RECT 74.460 32.870 74.830 33.180 ;
        RECT 77.710 32.960 78.030 33.270 ;
        RECT 78.620 32.960 78.940 33.270 ;
        RECT 81.810 33.180 82.100 33.420 ;
        RECT 80.210 32.870 80.580 33.180 ;
        RECT 83.460 32.960 83.780 33.270 ;
        RECT 84.370 32.960 84.690 33.270 ;
        RECT 87.560 33.180 87.850 33.420 ;
        RECT 85.960 32.870 86.330 33.180 ;
        RECT 89.210 32.960 89.530 33.270 ;
        RECT 90.120 32.960 90.440 33.270 ;
        RECT 93.310 33.180 93.600 33.420 ;
        RECT 91.710 32.870 92.080 33.180 ;
        RECT 3.360 31.370 3.650 31.630 ;
        RECT 1.260 31.150 1.580 31.210 ;
        RECT 3.430 31.150 3.570 31.370 ;
        RECT 4.930 31.290 5.250 31.600 ;
        RECT 6.570 31.290 6.890 31.600 ;
        RECT 7.480 31.290 7.800 31.600 ;
        RECT 9.110 31.370 9.400 31.630 ;
        RECT 9.180 31.150 9.320 31.370 ;
        RECT 10.680 31.290 11.000 31.600 ;
        RECT 12.320 31.290 12.640 31.600 ;
        RECT 13.230 31.290 13.550 31.600 ;
        RECT 14.860 31.370 15.150 31.630 ;
        RECT 14.930 31.150 15.070 31.370 ;
        RECT 16.430 31.290 16.750 31.600 ;
        RECT 18.070 31.290 18.390 31.600 ;
        RECT 18.980 31.290 19.300 31.600 ;
        RECT 20.610 31.370 20.900 31.630 ;
        RECT 20.680 31.150 20.820 31.370 ;
        RECT 22.180 31.290 22.500 31.600 ;
        RECT 23.820 31.290 24.140 31.600 ;
        RECT 24.730 31.290 25.050 31.600 ;
        RECT 26.360 31.370 26.650 31.630 ;
        RECT 26.430 31.150 26.570 31.370 ;
        RECT 27.930 31.290 28.250 31.600 ;
        RECT 29.570 31.290 29.890 31.600 ;
        RECT 30.480 31.290 30.800 31.600 ;
        RECT 32.110 31.370 32.400 31.630 ;
        RECT 32.180 31.150 32.320 31.370 ;
        RECT 33.680 31.290 34.000 31.600 ;
        RECT 35.320 31.290 35.640 31.600 ;
        RECT 36.230 31.290 36.550 31.600 ;
        RECT 37.860 31.370 38.150 31.630 ;
        RECT 37.930 31.150 38.070 31.370 ;
        RECT 39.430 31.290 39.750 31.600 ;
        RECT 41.070 31.290 41.390 31.600 ;
        RECT 41.980 31.290 42.300 31.600 ;
        RECT 43.610 31.370 43.900 31.630 ;
        RECT 43.680 31.150 43.820 31.370 ;
        RECT 45.180 31.290 45.500 31.600 ;
        RECT 46.820 31.290 47.140 31.600 ;
        RECT 47.730 31.290 48.050 31.600 ;
        RECT 49.360 31.370 49.650 31.630 ;
        RECT 49.430 31.150 49.570 31.370 ;
        RECT 50.930 31.290 51.250 31.600 ;
        RECT 52.570 31.290 52.890 31.600 ;
        RECT 53.480 31.290 53.800 31.600 ;
        RECT 55.110 31.370 55.400 31.630 ;
        RECT 55.180 31.150 55.320 31.370 ;
        RECT 56.680 31.290 57.000 31.600 ;
        RECT 58.320 31.290 58.640 31.600 ;
        RECT 59.230 31.290 59.550 31.600 ;
        RECT 60.860 31.370 61.150 31.630 ;
        RECT 60.930 31.150 61.070 31.370 ;
        RECT 62.430 31.290 62.750 31.600 ;
        RECT 64.070 31.290 64.390 31.600 ;
        RECT 64.980 31.290 65.300 31.600 ;
        RECT 66.610 31.370 66.900 31.630 ;
        RECT 66.680 31.150 66.820 31.370 ;
        RECT 68.180 31.290 68.500 31.600 ;
        RECT 69.820 31.290 70.140 31.600 ;
        RECT 70.730 31.290 71.050 31.600 ;
        RECT 72.360 31.370 72.650 31.630 ;
        RECT 72.430 31.150 72.570 31.370 ;
        RECT 73.930 31.290 74.250 31.600 ;
        RECT 75.570 31.290 75.890 31.600 ;
        RECT 76.480 31.290 76.800 31.600 ;
        RECT 78.110 31.370 78.400 31.630 ;
        RECT 78.180 31.150 78.320 31.370 ;
        RECT 79.680 31.290 80.000 31.600 ;
        RECT 81.320 31.290 81.640 31.600 ;
        RECT 82.230 31.290 82.550 31.600 ;
        RECT 83.860 31.370 84.150 31.630 ;
        RECT 83.930 31.150 84.070 31.370 ;
        RECT 85.430 31.290 85.750 31.600 ;
        RECT 87.070 31.290 87.390 31.600 ;
        RECT 87.980 31.290 88.300 31.600 ;
        RECT 89.610 31.370 89.900 31.630 ;
        RECT 89.680 31.150 89.820 31.370 ;
        RECT 91.180 31.290 91.500 31.600 ;
        RECT 92.820 31.290 93.140 31.600 ;
        RECT 93.730 31.290 94.050 31.600 ;
        RECT 1.260 31.010 94.660 31.150 ;
        RECT 1.260 30.950 1.580 31.010 ;
        RECT 2.960 30.550 3.280 30.860 ;
        RECT 3.870 30.550 4.190 30.860 ;
        RECT 7.060 30.770 7.350 31.010 ;
        RECT 5.460 30.460 5.830 30.770 ;
        RECT 8.710 30.550 9.030 30.860 ;
        RECT 9.620 30.550 9.940 30.860 ;
        RECT 12.810 30.770 13.100 31.010 ;
        RECT 11.210 30.460 11.580 30.770 ;
        RECT 14.460 30.550 14.780 30.860 ;
        RECT 15.370 30.550 15.690 30.860 ;
        RECT 18.560 30.770 18.850 31.010 ;
        RECT 16.960 30.460 17.330 30.770 ;
        RECT 20.210 30.550 20.530 30.860 ;
        RECT 21.120 30.550 21.440 30.860 ;
        RECT 24.310 30.770 24.600 31.010 ;
        RECT 22.710 30.460 23.080 30.770 ;
        RECT 25.960 30.550 26.280 30.860 ;
        RECT 26.870 30.550 27.190 30.860 ;
        RECT 30.060 30.770 30.350 31.010 ;
        RECT 28.460 30.460 28.830 30.770 ;
        RECT 31.710 30.550 32.030 30.860 ;
        RECT 32.620 30.550 32.940 30.860 ;
        RECT 35.810 30.770 36.100 31.010 ;
        RECT 34.210 30.460 34.580 30.770 ;
        RECT 37.460 30.550 37.780 30.860 ;
        RECT 38.370 30.550 38.690 30.860 ;
        RECT 41.560 30.770 41.850 31.010 ;
        RECT 39.960 30.460 40.330 30.770 ;
        RECT 43.210 30.550 43.530 30.860 ;
        RECT 44.120 30.550 44.440 30.860 ;
        RECT 47.310 30.770 47.600 31.010 ;
        RECT 45.710 30.460 46.080 30.770 ;
        RECT 48.960 30.550 49.280 30.860 ;
        RECT 49.870 30.550 50.190 30.860 ;
        RECT 53.060 30.770 53.350 31.010 ;
        RECT 51.460 30.460 51.830 30.770 ;
        RECT 54.710 30.550 55.030 30.860 ;
        RECT 55.620 30.550 55.940 30.860 ;
        RECT 58.810 30.770 59.100 31.010 ;
        RECT 57.210 30.460 57.580 30.770 ;
        RECT 60.460 30.550 60.780 30.860 ;
        RECT 61.370 30.550 61.690 30.860 ;
        RECT 64.560 30.770 64.850 31.010 ;
        RECT 62.960 30.460 63.330 30.770 ;
        RECT 66.210 30.550 66.530 30.860 ;
        RECT 67.120 30.550 67.440 30.860 ;
        RECT 70.310 30.770 70.600 31.010 ;
        RECT 68.710 30.460 69.080 30.770 ;
        RECT 71.960 30.550 72.280 30.860 ;
        RECT 72.870 30.550 73.190 30.860 ;
        RECT 76.060 30.770 76.350 31.010 ;
        RECT 74.460 30.460 74.830 30.770 ;
        RECT 77.710 30.550 78.030 30.860 ;
        RECT 78.620 30.550 78.940 30.860 ;
        RECT 81.810 30.770 82.100 31.010 ;
        RECT 80.210 30.460 80.580 30.770 ;
        RECT 83.460 30.550 83.780 30.860 ;
        RECT 84.370 30.550 84.690 30.860 ;
        RECT 87.560 30.770 87.850 31.010 ;
        RECT 85.960 30.460 86.330 30.770 ;
        RECT 89.210 30.550 89.530 30.860 ;
        RECT 90.120 30.550 90.440 30.860 ;
        RECT 93.310 30.770 93.600 31.010 ;
        RECT 91.710 30.460 92.080 30.770 ;
        RECT 3.360 28.960 3.650 29.220 ;
        RECT 1.260 28.740 1.580 28.800 ;
        RECT 3.430 28.740 3.570 28.960 ;
        RECT 4.930 28.880 5.250 29.190 ;
        RECT 6.570 28.880 6.890 29.190 ;
        RECT 7.480 28.880 7.800 29.190 ;
        RECT 9.110 28.960 9.400 29.220 ;
        RECT 9.180 28.740 9.320 28.960 ;
        RECT 10.680 28.880 11.000 29.190 ;
        RECT 12.320 28.880 12.640 29.190 ;
        RECT 13.230 28.880 13.550 29.190 ;
        RECT 14.860 28.960 15.150 29.220 ;
        RECT 14.930 28.740 15.070 28.960 ;
        RECT 16.430 28.880 16.750 29.190 ;
        RECT 18.070 28.880 18.390 29.190 ;
        RECT 18.980 28.880 19.300 29.190 ;
        RECT 20.610 28.960 20.900 29.220 ;
        RECT 20.680 28.740 20.820 28.960 ;
        RECT 22.180 28.880 22.500 29.190 ;
        RECT 23.820 28.880 24.140 29.190 ;
        RECT 24.730 28.880 25.050 29.190 ;
        RECT 26.360 28.960 26.650 29.220 ;
        RECT 26.430 28.740 26.570 28.960 ;
        RECT 27.930 28.880 28.250 29.190 ;
        RECT 29.570 28.880 29.890 29.190 ;
        RECT 30.480 28.880 30.800 29.190 ;
        RECT 32.110 28.960 32.400 29.220 ;
        RECT 32.180 28.740 32.320 28.960 ;
        RECT 33.680 28.880 34.000 29.190 ;
        RECT 35.320 28.880 35.640 29.190 ;
        RECT 36.230 28.880 36.550 29.190 ;
        RECT 37.860 28.960 38.150 29.220 ;
        RECT 37.930 28.740 38.070 28.960 ;
        RECT 39.430 28.880 39.750 29.190 ;
        RECT 41.070 28.880 41.390 29.190 ;
        RECT 41.980 28.880 42.300 29.190 ;
        RECT 43.610 28.960 43.900 29.220 ;
        RECT 43.680 28.740 43.820 28.960 ;
        RECT 45.180 28.880 45.500 29.190 ;
        RECT 46.820 28.880 47.140 29.190 ;
        RECT 47.730 28.880 48.050 29.190 ;
        RECT 49.360 28.960 49.650 29.220 ;
        RECT 49.430 28.740 49.570 28.960 ;
        RECT 50.930 28.880 51.250 29.190 ;
        RECT 52.570 28.880 52.890 29.190 ;
        RECT 53.480 28.880 53.800 29.190 ;
        RECT 55.110 28.960 55.400 29.220 ;
        RECT 55.180 28.740 55.320 28.960 ;
        RECT 56.680 28.880 57.000 29.190 ;
        RECT 58.320 28.880 58.640 29.190 ;
        RECT 59.230 28.880 59.550 29.190 ;
        RECT 60.860 28.960 61.150 29.220 ;
        RECT 60.930 28.740 61.070 28.960 ;
        RECT 62.430 28.880 62.750 29.190 ;
        RECT 64.070 28.880 64.390 29.190 ;
        RECT 64.980 28.880 65.300 29.190 ;
        RECT 66.610 28.960 66.900 29.220 ;
        RECT 66.680 28.740 66.820 28.960 ;
        RECT 68.180 28.880 68.500 29.190 ;
        RECT 69.820 28.880 70.140 29.190 ;
        RECT 70.730 28.880 71.050 29.190 ;
        RECT 72.360 28.960 72.650 29.220 ;
        RECT 72.430 28.740 72.570 28.960 ;
        RECT 73.930 28.880 74.250 29.190 ;
        RECT 75.570 28.880 75.890 29.190 ;
        RECT 76.480 28.880 76.800 29.190 ;
        RECT 78.110 28.960 78.400 29.220 ;
        RECT 78.180 28.740 78.320 28.960 ;
        RECT 79.680 28.880 80.000 29.190 ;
        RECT 81.320 28.880 81.640 29.190 ;
        RECT 82.230 28.880 82.550 29.190 ;
        RECT 83.860 28.960 84.150 29.220 ;
        RECT 83.930 28.740 84.070 28.960 ;
        RECT 85.430 28.880 85.750 29.190 ;
        RECT 87.070 28.880 87.390 29.190 ;
        RECT 87.980 28.880 88.300 29.190 ;
        RECT 89.610 28.960 89.900 29.220 ;
        RECT 89.680 28.740 89.820 28.960 ;
        RECT 91.180 28.880 91.500 29.190 ;
        RECT 92.820 28.880 93.140 29.190 ;
        RECT 93.730 28.880 94.050 29.190 ;
        RECT 1.260 28.600 94.660 28.740 ;
        RECT 1.260 28.540 1.580 28.600 ;
        RECT 7.140 28.310 7.280 28.600 ;
        RECT 12.890 28.310 13.030 28.600 ;
        RECT 18.640 28.310 18.780 28.600 ;
        RECT 24.390 28.310 24.530 28.600 ;
        RECT 30.140 28.310 30.280 28.600 ;
        RECT 35.890 28.310 36.030 28.600 ;
        RECT 41.640 28.310 41.780 28.600 ;
        RECT 47.390 28.310 47.530 28.600 ;
        RECT 53.140 28.310 53.280 28.600 ;
        RECT 58.890 28.310 59.030 28.600 ;
        RECT 64.640 28.310 64.780 28.600 ;
        RECT 70.390 28.310 70.530 28.600 ;
        RECT 76.140 28.310 76.280 28.600 ;
        RECT 81.890 28.310 82.030 28.600 ;
        RECT 87.640 28.310 87.780 28.600 ;
        RECT 93.390 28.310 93.530 28.600 ;
        RECT 7.060 28.060 7.350 28.310 ;
        RECT 12.810 28.060 13.100 28.310 ;
        RECT 18.560 28.060 18.850 28.310 ;
        RECT 24.310 28.060 24.600 28.310 ;
        RECT 30.060 28.060 30.350 28.310 ;
        RECT 35.810 28.060 36.100 28.310 ;
        RECT 41.560 28.060 41.850 28.310 ;
        RECT 47.310 28.060 47.600 28.310 ;
        RECT 53.060 28.060 53.350 28.310 ;
        RECT 58.810 28.060 59.100 28.310 ;
        RECT 64.560 28.060 64.850 28.310 ;
        RECT 70.310 28.060 70.600 28.310 ;
        RECT 76.060 28.060 76.350 28.310 ;
        RECT 81.810 28.060 82.100 28.310 ;
        RECT 87.560 28.060 87.850 28.310 ;
        RECT 93.310 28.060 93.600 28.310 ;
        RECT 2.960 27.740 3.280 28.050 ;
        RECT 3.870 27.740 4.190 28.050 ;
        RECT 5.460 27.650 5.830 27.960 ;
        RECT 8.710 27.740 9.030 28.050 ;
        RECT 9.620 27.740 9.940 28.050 ;
        RECT 11.210 27.650 11.580 27.960 ;
        RECT 14.460 27.740 14.780 28.050 ;
        RECT 15.370 27.740 15.690 28.050 ;
        RECT 16.960 27.650 17.330 27.960 ;
        RECT 20.210 27.740 20.530 28.050 ;
        RECT 21.120 27.740 21.440 28.050 ;
        RECT 22.710 27.650 23.080 27.960 ;
        RECT 25.960 27.740 26.280 28.050 ;
        RECT 26.870 27.740 27.190 28.050 ;
        RECT 28.460 27.650 28.830 27.960 ;
        RECT 31.710 27.740 32.030 28.050 ;
        RECT 32.620 27.740 32.940 28.050 ;
        RECT 34.210 27.650 34.580 27.960 ;
        RECT 37.460 27.740 37.780 28.050 ;
        RECT 38.370 27.740 38.690 28.050 ;
        RECT 39.960 27.650 40.330 27.960 ;
        RECT 43.210 27.740 43.530 28.050 ;
        RECT 44.120 27.740 44.440 28.050 ;
        RECT 45.710 27.650 46.080 27.960 ;
        RECT 48.960 27.740 49.280 28.050 ;
        RECT 49.870 27.740 50.190 28.050 ;
        RECT 51.460 27.650 51.830 27.960 ;
        RECT 54.710 27.740 55.030 28.050 ;
        RECT 55.620 27.740 55.940 28.050 ;
        RECT 57.210 27.650 57.580 27.960 ;
        RECT 60.460 27.740 60.780 28.050 ;
        RECT 61.370 27.740 61.690 28.050 ;
        RECT 62.960 27.650 63.330 27.960 ;
        RECT 66.210 27.740 66.530 28.050 ;
        RECT 67.120 27.740 67.440 28.050 ;
        RECT 68.710 27.650 69.080 27.960 ;
        RECT 71.960 27.740 72.280 28.050 ;
        RECT 72.870 27.740 73.190 28.050 ;
        RECT 74.460 27.650 74.830 27.960 ;
        RECT 77.710 27.740 78.030 28.050 ;
        RECT 78.620 27.740 78.940 28.050 ;
        RECT 80.210 27.650 80.580 27.960 ;
        RECT 83.460 27.740 83.780 28.050 ;
        RECT 84.370 27.740 84.690 28.050 ;
        RECT 85.960 27.650 86.330 27.960 ;
        RECT 89.210 27.740 89.530 28.050 ;
        RECT 90.120 27.740 90.440 28.050 ;
        RECT 91.710 27.650 92.080 27.960 ;
        RECT 3.360 26.150 3.650 26.410 ;
        RECT 1.250 25.930 1.570 25.990 ;
        RECT 3.430 25.930 3.570 26.150 ;
        RECT 4.930 26.070 5.250 26.380 ;
        RECT 6.570 26.070 6.890 26.380 ;
        RECT 7.480 26.070 7.800 26.380 ;
        RECT 9.110 26.150 9.400 26.410 ;
        RECT 9.180 25.930 9.320 26.150 ;
        RECT 10.680 26.070 11.000 26.380 ;
        RECT 12.320 26.070 12.640 26.380 ;
        RECT 13.230 26.070 13.550 26.380 ;
        RECT 14.860 26.150 15.150 26.410 ;
        RECT 14.930 25.930 15.070 26.150 ;
        RECT 16.430 26.070 16.750 26.380 ;
        RECT 18.070 26.070 18.390 26.380 ;
        RECT 18.980 26.070 19.300 26.380 ;
        RECT 20.610 26.150 20.900 26.410 ;
        RECT 20.680 25.930 20.820 26.150 ;
        RECT 22.180 26.070 22.500 26.380 ;
        RECT 23.820 26.070 24.140 26.380 ;
        RECT 24.730 26.070 25.050 26.380 ;
        RECT 26.360 26.150 26.650 26.410 ;
        RECT 26.430 25.930 26.570 26.150 ;
        RECT 27.930 26.070 28.250 26.380 ;
        RECT 29.570 26.070 29.890 26.380 ;
        RECT 30.480 26.070 30.800 26.380 ;
        RECT 32.110 26.150 32.400 26.410 ;
        RECT 32.180 25.930 32.320 26.150 ;
        RECT 33.680 26.070 34.000 26.380 ;
        RECT 35.320 26.070 35.640 26.380 ;
        RECT 36.230 26.070 36.550 26.380 ;
        RECT 37.860 26.150 38.150 26.410 ;
        RECT 37.930 25.930 38.070 26.150 ;
        RECT 39.430 26.070 39.750 26.380 ;
        RECT 41.070 26.070 41.390 26.380 ;
        RECT 41.980 26.070 42.300 26.380 ;
        RECT 43.610 26.150 43.900 26.410 ;
        RECT 43.680 25.930 43.820 26.150 ;
        RECT 45.180 26.070 45.500 26.380 ;
        RECT 46.820 26.070 47.140 26.380 ;
        RECT 47.730 26.070 48.050 26.380 ;
        RECT 49.360 26.150 49.650 26.410 ;
        RECT 49.430 25.930 49.570 26.150 ;
        RECT 50.930 26.070 51.250 26.380 ;
        RECT 52.570 26.070 52.890 26.380 ;
        RECT 53.480 26.070 53.800 26.380 ;
        RECT 55.110 26.150 55.400 26.410 ;
        RECT 55.180 25.930 55.320 26.150 ;
        RECT 56.680 26.070 57.000 26.380 ;
        RECT 58.320 26.070 58.640 26.380 ;
        RECT 59.230 26.070 59.550 26.380 ;
        RECT 60.860 26.150 61.150 26.410 ;
        RECT 60.930 25.930 61.070 26.150 ;
        RECT 62.430 26.070 62.750 26.380 ;
        RECT 64.070 26.070 64.390 26.380 ;
        RECT 64.980 26.070 65.300 26.380 ;
        RECT 66.610 26.150 66.900 26.410 ;
        RECT 66.680 25.930 66.820 26.150 ;
        RECT 68.180 26.070 68.500 26.380 ;
        RECT 69.820 26.070 70.140 26.380 ;
        RECT 70.730 26.070 71.050 26.380 ;
        RECT 72.360 26.150 72.650 26.410 ;
        RECT 72.430 25.930 72.570 26.150 ;
        RECT 73.930 26.070 74.250 26.380 ;
        RECT 75.570 26.070 75.890 26.380 ;
        RECT 76.480 26.070 76.800 26.380 ;
        RECT 78.110 26.150 78.400 26.410 ;
        RECT 78.180 25.930 78.320 26.150 ;
        RECT 79.680 26.070 80.000 26.380 ;
        RECT 81.320 26.070 81.640 26.380 ;
        RECT 82.230 26.070 82.550 26.380 ;
        RECT 83.860 26.150 84.150 26.410 ;
        RECT 83.930 25.930 84.070 26.150 ;
        RECT 85.430 26.070 85.750 26.380 ;
        RECT 87.070 26.070 87.390 26.380 ;
        RECT 87.980 26.070 88.300 26.380 ;
        RECT 89.610 26.150 89.900 26.410 ;
        RECT 89.680 25.930 89.820 26.150 ;
        RECT 91.180 26.070 91.500 26.380 ;
        RECT 92.820 26.070 93.140 26.380 ;
        RECT 93.730 26.070 94.050 26.380 ;
        RECT 1.250 25.790 94.660 25.930 ;
        RECT 1.250 25.730 1.570 25.790 ;
        RECT 2.960 25.330 3.280 25.640 ;
        RECT 3.870 25.330 4.190 25.640 ;
        RECT 7.060 25.550 7.350 25.790 ;
        RECT 5.460 25.240 5.830 25.550 ;
        RECT 8.710 25.330 9.030 25.640 ;
        RECT 9.620 25.330 9.940 25.640 ;
        RECT 12.810 25.550 13.100 25.790 ;
        RECT 11.210 25.240 11.580 25.550 ;
        RECT 14.460 25.330 14.780 25.640 ;
        RECT 15.370 25.330 15.690 25.640 ;
        RECT 18.560 25.550 18.850 25.790 ;
        RECT 16.960 25.240 17.330 25.550 ;
        RECT 20.210 25.330 20.530 25.640 ;
        RECT 21.120 25.330 21.440 25.640 ;
        RECT 24.310 25.550 24.600 25.790 ;
        RECT 22.710 25.240 23.080 25.550 ;
        RECT 25.960 25.330 26.280 25.640 ;
        RECT 26.870 25.330 27.190 25.640 ;
        RECT 30.060 25.550 30.350 25.790 ;
        RECT 28.460 25.240 28.830 25.550 ;
        RECT 31.710 25.330 32.030 25.640 ;
        RECT 32.620 25.330 32.940 25.640 ;
        RECT 35.810 25.550 36.100 25.790 ;
        RECT 34.210 25.240 34.580 25.550 ;
        RECT 37.460 25.330 37.780 25.640 ;
        RECT 38.370 25.330 38.690 25.640 ;
        RECT 41.560 25.550 41.850 25.790 ;
        RECT 39.960 25.240 40.330 25.550 ;
        RECT 43.210 25.330 43.530 25.640 ;
        RECT 44.120 25.330 44.440 25.640 ;
        RECT 47.310 25.550 47.600 25.790 ;
        RECT 45.710 25.240 46.080 25.550 ;
        RECT 48.960 25.330 49.280 25.640 ;
        RECT 49.870 25.330 50.190 25.640 ;
        RECT 53.060 25.550 53.350 25.790 ;
        RECT 51.460 25.240 51.830 25.550 ;
        RECT 54.710 25.330 55.030 25.640 ;
        RECT 55.620 25.330 55.940 25.640 ;
        RECT 58.810 25.550 59.100 25.790 ;
        RECT 57.210 25.240 57.580 25.550 ;
        RECT 60.460 25.330 60.780 25.640 ;
        RECT 61.370 25.330 61.690 25.640 ;
        RECT 64.560 25.550 64.850 25.790 ;
        RECT 62.960 25.240 63.330 25.550 ;
        RECT 66.210 25.330 66.530 25.640 ;
        RECT 67.120 25.330 67.440 25.640 ;
        RECT 70.310 25.550 70.600 25.790 ;
        RECT 68.710 25.240 69.080 25.550 ;
        RECT 71.960 25.330 72.280 25.640 ;
        RECT 72.870 25.330 73.190 25.640 ;
        RECT 76.060 25.550 76.350 25.790 ;
        RECT 74.460 25.240 74.830 25.550 ;
        RECT 77.710 25.330 78.030 25.640 ;
        RECT 78.620 25.330 78.940 25.640 ;
        RECT 81.810 25.550 82.100 25.790 ;
        RECT 80.210 25.240 80.580 25.550 ;
        RECT 83.460 25.330 83.780 25.640 ;
        RECT 84.370 25.330 84.690 25.640 ;
        RECT 87.560 25.550 87.850 25.790 ;
        RECT 85.960 25.240 86.330 25.550 ;
        RECT 89.210 25.330 89.530 25.640 ;
        RECT 90.120 25.330 90.440 25.640 ;
        RECT 93.310 25.550 93.600 25.790 ;
        RECT 91.710 25.240 92.080 25.550 ;
        RECT 3.360 23.740 3.650 24.000 ;
        RECT 1.260 23.520 1.580 23.580 ;
        RECT 3.430 23.520 3.570 23.740 ;
        RECT 4.930 23.660 5.250 23.970 ;
        RECT 6.570 23.660 6.890 23.970 ;
        RECT 7.480 23.660 7.800 23.970 ;
        RECT 9.110 23.740 9.400 24.000 ;
        RECT 9.180 23.520 9.320 23.740 ;
        RECT 10.680 23.660 11.000 23.970 ;
        RECT 12.320 23.660 12.640 23.970 ;
        RECT 13.230 23.660 13.550 23.970 ;
        RECT 14.860 23.740 15.150 24.000 ;
        RECT 14.930 23.520 15.070 23.740 ;
        RECT 16.430 23.660 16.750 23.970 ;
        RECT 18.070 23.660 18.390 23.970 ;
        RECT 18.980 23.660 19.300 23.970 ;
        RECT 20.610 23.740 20.900 24.000 ;
        RECT 20.680 23.520 20.820 23.740 ;
        RECT 22.180 23.660 22.500 23.970 ;
        RECT 23.820 23.660 24.140 23.970 ;
        RECT 24.730 23.660 25.050 23.970 ;
        RECT 26.360 23.740 26.650 24.000 ;
        RECT 26.430 23.520 26.570 23.740 ;
        RECT 27.930 23.660 28.250 23.970 ;
        RECT 29.570 23.660 29.890 23.970 ;
        RECT 30.480 23.660 30.800 23.970 ;
        RECT 32.110 23.740 32.400 24.000 ;
        RECT 32.180 23.520 32.320 23.740 ;
        RECT 33.680 23.660 34.000 23.970 ;
        RECT 35.320 23.660 35.640 23.970 ;
        RECT 36.230 23.660 36.550 23.970 ;
        RECT 37.860 23.740 38.150 24.000 ;
        RECT 37.930 23.520 38.070 23.740 ;
        RECT 39.430 23.660 39.750 23.970 ;
        RECT 41.070 23.660 41.390 23.970 ;
        RECT 41.980 23.660 42.300 23.970 ;
        RECT 43.610 23.740 43.900 24.000 ;
        RECT 43.680 23.520 43.820 23.740 ;
        RECT 45.180 23.660 45.500 23.970 ;
        RECT 46.820 23.660 47.140 23.970 ;
        RECT 47.730 23.660 48.050 23.970 ;
        RECT 49.360 23.740 49.650 24.000 ;
        RECT 49.430 23.520 49.570 23.740 ;
        RECT 50.930 23.660 51.250 23.970 ;
        RECT 52.570 23.660 52.890 23.970 ;
        RECT 53.480 23.660 53.800 23.970 ;
        RECT 55.110 23.740 55.400 24.000 ;
        RECT 55.180 23.520 55.320 23.740 ;
        RECT 56.680 23.660 57.000 23.970 ;
        RECT 58.320 23.660 58.640 23.970 ;
        RECT 59.230 23.660 59.550 23.970 ;
        RECT 60.860 23.740 61.150 24.000 ;
        RECT 60.930 23.520 61.070 23.740 ;
        RECT 62.430 23.660 62.750 23.970 ;
        RECT 64.070 23.660 64.390 23.970 ;
        RECT 64.980 23.660 65.300 23.970 ;
        RECT 66.610 23.740 66.900 24.000 ;
        RECT 66.680 23.520 66.820 23.740 ;
        RECT 68.180 23.660 68.500 23.970 ;
        RECT 69.820 23.660 70.140 23.970 ;
        RECT 70.730 23.660 71.050 23.970 ;
        RECT 72.360 23.740 72.650 24.000 ;
        RECT 72.430 23.520 72.570 23.740 ;
        RECT 73.930 23.660 74.250 23.970 ;
        RECT 75.570 23.660 75.890 23.970 ;
        RECT 76.480 23.660 76.800 23.970 ;
        RECT 78.110 23.740 78.400 24.000 ;
        RECT 78.180 23.520 78.320 23.740 ;
        RECT 79.680 23.660 80.000 23.970 ;
        RECT 81.320 23.660 81.640 23.970 ;
        RECT 82.230 23.660 82.550 23.970 ;
        RECT 83.860 23.740 84.150 24.000 ;
        RECT 83.930 23.520 84.070 23.740 ;
        RECT 85.430 23.660 85.750 23.970 ;
        RECT 87.070 23.660 87.390 23.970 ;
        RECT 87.980 23.660 88.300 23.970 ;
        RECT 89.610 23.740 89.900 24.000 ;
        RECT 89.680 23.520 89.820 23.740 ;
        RECT 91.180 23.660 91.500 23.970 ;
        RECT 92.820 23.660 93.140 23.970 ;
        RECT 93.730 23.660 94.050 23.970 ;
        RECT 1.260 23.380 94.660 23.520 ;
        RECT 1.260 23.320 1.580 23.380 ;
        RECT 2.960 22.920 3.280 23.230 ;
        RECT 3.870 22.920 4.190 23.230 ;
        RECT 7.060 23.140 7.350 23.380 ;
        RECT 5.460 22.830 5.830 23.140 ;
        RECT 8.710 22.920 9.030 23.230 ;
        RECT 9.620 22.920 9.940 23.230 ;
        RECT 12.810 23.140 13.100 23.380 ;
        RECT 11.210 22.830 11.580 23.140 ;
        RECT 14.460 22.920 14.780 23.230 ;
        RECT 15.370 22.920 15.690 23.230 ;
        RECT 18.560 23.140 18.850 23.380 ;
        RECT 16.960 22.830 17.330 23.140 ;
        RECT 20.210 22.920 20.530 23.230 ;
        RECT 21.120 22.920 21.440 23.230 ;
        RECT 24.310 23.140 24.600 23.380 ;
        RECT 22.710 22.830 23.080 23.140 ;
        RECT 25.960 22.920 26.280 23.230 ;
        RECT 26.870 22.920 27.190 23.230 ;
        RECT 30.060 23.140 30.350 23.380 ;
        RECT 28.460 22.830 28.830 23.140 ;
        RECT 31.710 22.920 32.030 23.230 ;
        RECT 32.620 22.920 32.940 23.230 ;
        RECT 35.810 23.140 36.100 23.380 ;
        RECT 34.210 22.830 34.580 23.140 ;
        RECT 37.460 22.920 37.780 23.230 ;
        RECT 38.370 22.920 38.690 23.230 ;
        RECT 41.560 23.140 41.850 23.380 ;
        RECT 39.960 22.830 40.330 23.140 ;
        RECT 43.210 22.920 43.530 23.230 ;
        RECT 44.120 22.920 44.440 23.230 ;
        RECT 47.310 23.140 47.600 23.380 ;
        RECT 45.710 22.830 46.080 23.140 ;
        RECT 48.960 22.920 49.280 23.230 ;
        RECT 49.870 22.920 50.190 23.230 ;
        RECT 53.060 23.140 53.350 23.380 ;
        RECT 51.460 22.830 51.830 23.140 ;
        RECT 54.710 22.920 55.030 23.230 ;
        RECT 55.620 22.920 55.940 23.230 ;
        RECT 58.810 23.140 59.100 23.380 ;
        RECT 57.210 22.830 57.580 23.140 ;
        RECT 60.460 22.920 60.780 23.230 ;
        RECT 61.370 22.920 61.690 23.230 ;
        RECT 64.560 23.140 64.850 23.380 ;
        RECT 62.960 22.830 63.330 23.140 ;
        RECT 66.210 22.920 66.530 23.230 ;
        RECT 67.120 22.920 67.440 23.230 ;
        RECT 70.310 23.140 70.600 23.380 ;
        RECT 68.710 22.830 69.080 23.140 ;
        RECT 71.960 22.920 72.280 23.230 ;
        RECT 72.870 22.920 73.190 23.230 ;
        RECT 76.060 23.140 76.350 23.380 ;
        RECT 74.460 22.830 74.830 23.140 ;
        RECT 77.710 22.920 78.030 23.230 ;
        RECT 78.620 22.920 78.940 23.230 ;
        RECT 81.810 23.140 82.100 23.380 ;
        RECT 80.210 22.830 80.580 23.140 ;
        RECT 83.460 22.920 83.780 23.230 ;
        RECT 84.370 22.920 84.690 23.230 ;
        RECT 87.560 23.140 87.850 23.380 ;
        RECT 85.960 22.830 86.330 23.140 ;
        RECT 89.210 22.920 89.530 23.230 ;
        RECT 90.120 22.920 90.440 23.230 ;
        RECT 93.310 23.140 93.600 23.380 ;
        RECT 91.710 22.830 92.080 23.140 ;
        RECT 3.360 21.330 3.650 21.590 ;
        RECT 1.260 21.110 1.580 21.170 ;
        RECT 3.430 21.110 3.570 21.330 ;
        RECT 4.930 21.250 5.250 21.560 ;
        RECT 6.570 21.250 6.890 21.560 ;
        RECT 7.480 21.250 7.800 21.560 ;
        RECT 9.110 21.330 9.400 21.590 ;
        RECT 9.180 21.110 9.320 21.330 ;
        RECT 10.680 21.250 11.000 21.560 ;
        RECT 12.320 21.250 12.640 21.560 ;
        RECT 13.230 21.250 13.550 21.560 ;
        RECT 14.860 21.330 15.150 21.590 ;
        RECT 14.930 21.110 15.070 21.330 ;
        RECT 16.430 21.250 16.750 21.560 ;
        RECT 18.070 21.250 18.390 21.560 ;
        RECT 18.980 21.250 19.300 21.560 ;
        RECT 20.610 21.330 20.900 21.590 ;
        RECT 20.680 21.110 20.820 21.330 ;
        RECT 22.180 21.250 22.500 21.560 ;
        RECT 23.820 21.250 24.140 21.560 ;
        RECT 24.730 21.250 25.050 21.560 ;
        RECT 26.360 21.330 26.650 21.590 ;
        RECT 26.430 21.110 26.570 21.330 ;
        RECT 27.930 21.250 28.250 21.560 ;
        RECT 29.570 21.250 29.890 21.560 ;
        RECT 30.480 21.250 30.800 21.560 ;
        RECT 32.110 21.330 32.400 21.590 ;
        RECT 32.180 21.110 32.320 21.330 ;
        RECT 33.680 21.250 34.000 21.560 ;
        RECT 35.320 21.250 35.640 21.560 ;
        RECT 36.230 21.250 36.550 21.560 ;
        RECT 37.860 21.330 38.150 21.590 ;
        RECT 37.930 21.110 38.070 21.330 ;
        RECT 39.430 21.250 39.750 21.560 ;
        RECT 41.070 21.250 41.390 21.560 ;
        RECT 41.980 21.250 42.300 21.560 ;
        RECT 43.610 21.330 43.900 21.590 ;
        RECT 43.680 21.110 43.820 21.330 ;
        RECT 45.180 21.250 45.500 21.560 ;
        RECT 46.820 21.250 47.140 21.560 ;
        RECT 47.730 21.250 48.050 21.560 ;
        RECT 49.360 21.330 49.650 21.590 ;
        RECT 49.430 21.110 49.570 21.330 ;
        RECT 50.930 21.250 51.250 21.560 ;
        RECT 52.570 21.250 52.890 21.560 ;
        RECT 53.480 21.250 53.800 21.560 ;
        RECT 55.110 21.330 55.400 21.590 ;
        RECT 55.180 21.110 55.320 21.330 ;
        RECT 56.680 21.250 57.000 21.560 ;
        RECT 58.320 21.250 58.640 21.560 ;
        RECT 59.230 21.250 59.550 21.560 ;
        RECT 60.860 21.330 61.150 21.590 ;
        RECT 60.930 21.110 61.070 21.330 ;
        RECT 62.430 21.250 62.750 21.560 ;
        RECT 64.070 21.250 64.390 21.560 ;
        RECT 64.980 21.250 65.300 21.560 ;
        RECT 66.610 21.330 66.900 21.590 ;
        RECT 66.680 21.110 66.820 21.330 ;
        RECT 68.180 21.250 68.500 21.560 ;
        RECT 69.820 21.250 70.140 21.560 ;
        RECT 70.730 21.250 71.050 21.560 ;
        RECT 72.360 21.330 72.650 21.590 ;
        RECT 72.430 21.110 72.570 21.330 ;
        RECT 73.930 21.250 74.250 21.560 ;
        RECT 75.570 21.250 75.890 21.560 ;
        RECT 76.480 21.250 76.800 21.560 ;
        RECT 78.110 21.330 78.400 21.590 ;
        RECT 78.180 21.110 78.320 21.330 ;
        RECT 79.680 21.250 80.000 21.560 ;
        RECT 81.320 21.250 81.640 21.560 ;
        RECT 82.230 21.250 82.550 21.560 ;
        RECT 83.860 21.330 84.150 21.590 ;
        RECT 83.930 21.110 84.070 21.330 ;
        RECT 85.430 21.250 85.750 21.560 ;
        RECT 87.070 21.250 87.390 21.560 ;
        RECT 87.980 21.250 88.300 21.560 ;
        RECT 89.610 21.330 89.900 21.590 ;
        RECT 89.680 21.110 89.820 21.330 ;
        RECT 91.180 21.250 91.500 21.560 ;
        RECT 92.820 21.250 93.140 21.560 ;
        RECT 93.730 21.250 94.050 21.560 ;
        RECT 1.260 20.970 94.660 21.110 ;
        RECT 1.260 20.910 1.580 20.970 ;
        RECT 2.960 20.510 3.280 20.820 ;
        RECT 3.870 20.510 4.190 20.820 ;
        RECT 7.060 20.730 7.350 20.970 ;
        RECT 5.460 20.420 5.830 20.730 ;
        RECT 8.710 20.510 9.030 20.820 ;
        RECT 9.620 20.510 9.940 20.820 ;
        RECT 12.810 20.730 13.100 20.970 ;
        RECT 11.210 20.420 11.580 20.730 ;
        RECT 14.460 20.510 14.780 20.820 ;
        RECT 15.370 20.510 15.690 20.820 ;
        RECT 18.560 20.730 18.850 20.970 ;
        RECT 16.960 20.420 17.330 20.730 ;
        RECT 20.210 20.510 20.530 20.820 ;
        RECT 21.120 20.510 21.440 20.820 ;
        RECT 24.310 20.730 24.600 20.970 ;
        RECT 22.710 20.420 23.080 20.730 ;
        RECT 25.960 20.510 26.280 20.820 ;
        RECT 26.870 20.510 27.190 20.820 ;
        RECT 30.060 20.730 30.350 20.970 ;
        RECT 28.460 20.420 28.830 20.730 ;
        RECT 31.710 20.510 32.030 20.820 ;
        RECT 32.620 20.510 32.940 20.820 ;
        RECT 35.810 20.730 36.100 20.970 ;
        RECT 34.210 20.420 34.580 20.730 ;
        RECT 37.460 20.510 37.780 20.820 ;
        RECT 38.370 20.510 38.690 20.820 ;
        RECT 41.560 20.730 41.850 20.970 ;
        RECT 39.960 20.420 40.330 20.730 ;
        RECT 43.210 20.510 43.530 20.820 ;
        RECT 44.120 20.510 44.440 20.820 ;
        RECT 47.310 20.730 47.600 20.970 ;
        RECT 45.710 20.420 46.080 20.730 ;
        RECT 48.960 20.510 49.280 20.820 ;
        RECT 49.870 20.510 50.190 20.820 ;
        RECT 53.060 20.730 53.350 20.970 ;
        RECT 51.460 20.420 51.830 20.730 ;
        RECT 54.710 20.510 55.030 20.820 ;
        RECT 55.620 20.510 55.940 20.820 ;
        RECT 58.810 20.730 59.100 20.970 ;
        RECT 57.210 20.420 57.580 20.730 ;
        RECT 60.460 20.510 60.780 20.820 ;
        RECT 61.370 20.510 61.690 20.820 ;
        RECT 64.560 20.730 64.850 20.970 ;
        RECT 62.960 20.420 63.330 20.730 ;
        RECT 66.210 20.510 66.530 20.820 ;
        RECT 67.120 20.510 67.440 20.820 ;
        RECT 70.310 20.730 70.600 20.970 ;
        RECT 68.710 20.420 69.080 20.730 ;
        RECT 71.960 20.510 72.280 20.820 ;
        RECT 72.870 20.510 73.190 20.820 ;
        RECT 76.060 20.730 76.350 20.970 ;
        RECT 74.460 20.420 74.830 20.730 ;
        RECT 77.710 20.510 78.030 20.820 ;
        RECT 78.620 20.510 78.940 20.820 ;
        RECT 81.810 20.730 82.100 20.970 ;
        RECT 80.210 20.420 80.580 20.730 ;
        RECT 83.460 20.510 83.780 20.820 ;
        RECT 84.370 20.510 84.690 20.820 ;
        RECT 87.560 20.730 87.850 20.970 ;
        RECT 85.960 20.420 86.330 20.730 ;
        RECT 89.210 20.510 89.530 20.820 ;
        RECT 90.120 20.510 90.440 20.820 ;
        RECT 93.310 20.730 93.600 20.970 ;
        RECT 91.710 20.420 92.080 20.730 ;
        RECT 3.360 18.920 3.650 19.180 ;
        RECT 1.260 18.700 1.580 18.760 ;
        RECT 3.430 18.700 3.570 18.920 ;
        RECT 4.930 18.840 5.250 19.150 ;
        RECT 6.570 18.840 6.890 19.150 ;
        RECT 7.480 18.840 7.800 19.150 ;
        RECT 9.110 18.920 9.400 19.180 ;
        RECT 9.180 18.700 9.320 18.920 ;
        RECT 10.680 18.840 11.000 19.150 ;
        RECT 12.320 18.840 12.640 19.150 ;
        RECT 13.230 18.840 13.550 19.150 ;
        RECT 14.860 18.920 15.150 19.180 ;
        RECT 14.930 18.700 15.070 18.920 ;
        RECT 16.430 18.840 16.750 19.150 ;
        RECT 18.070 18.840 18.390 19.150 ;
        RECT 18.980 18.840 19.300 19.150 ;
        RECT 20.610 18.920 20.900 19.180 ;
        RECT 20.680 18.700 20.820 18.920 ;
        RECT 22.180 18.840 22.500 19.150 ;
        RECT 23.820 18.840 24.140 19.150 ;
        RECT 24.730 18.840 25.050 19.150 ;
        RECT 26.360 18.920 26.650 19.180 ;
        RECT 26.430 18.700 26.570 18.920 ;
        RECT 27.930 18.840 28.250 19.150 ;
        RECT 29.570 18.840 29.890 19.150 ;
        RECT 30.480 18.840 30.800 19.150 ;
        RECT 32.110 18.920 32.400 19.180 ;
        RECT 32.180 18.700 32.320 18.920 ;
        RECT 33.680 18.840 34.000 19.150 ;
        RECT 35.320 18.840 35.640 19.150 ;
        RECT 36.230 18.840 36.550 19.150 ;
        RECT 37.860 18.920 38.150 19.180 ;
        RECT 37.930 18.700 38.070 18.920 ;
        RECT 39.430 18.840 39.750 19.150 ;
        RECT 41.070 18.840 41.390 19.150 ;
        RECT 41.980 18.840 42.300 19.150 ;
        RECT 43.610 18.920 43.900 19.180 ;
        RECT 43.680 18.700 43.820 18.920 ;
        RECT 45.180 18.840 45.500 19.150 ;
        RECT 46.820 18.840 47.140 19.150 ;
        RECT 47.730 18.840 48.050 19.150 ;
        RECT 49.360 18.920 49.650 19.180 ;
        RECT 49.430 18.700 49.570 18.920 ;
        RECT 50.930 18.840 51.250 19.150 ;
        RECT 52.570 18.840 52.890 19.150 ;
        RECT 53.480 18.840 53.800 19.150 ;
        RECT 55.110 18.920 55.400 19.180 ;
        RECT 55.180 18.700 55.320 18.920 ;
        RECT 56.680 18.840 57.000 19.150 ;
        RECT 58.320 18.840 58.640 19.150 ;
        RECT 59.230 18.840 59.550 19.150 ;
        RECT 60.860 18.920 61.150 19.180 ;
        RECT 60.930 18.700 61.070 18.920 ;
        RECT 62.430 18.840 62.750 19.150 ;
        RECT 64.070 18.840 64.390 19.150 ;
        RECT 64.980 18.840 65.300 19.150 ;
        RECT 66.610 18.920 66.900 19.180 ;
        RECT 66.680 18.700 66.820 18.920 ;
        RECT 68.180 18.840 68.500 19.150 ;
        RECT 69.820 18.840 70.140 19.150 ;
        RECT 70.730 18.840 71.050 19.150 ;
        RECT 72.360 18.920 72.650 19.180 ;
        RECT 72.430 18.700 72.570 18.920 ;
        RECT 73.930 18.840 74.250 19.150 ;
        RECT 75.570 18.840 75.890 19.150 ;
        RECT 76.480 18.840 76.800 19.150 ;
        RECT 78.110 18.920 78.400 19.180 ;
        RECT 78.180 18.700 78.320 18.920 ;
        RECT 79.680 18.840 80.000 19.150 ;
        RECT 81.320 18.840 81.640 19.150 ;
        RECT 82.230 18.840 82.550 19.150 ;
        RECT 83.860 18.920 84.150 19.180 ;
        RECT 83.930 18.700 84.070 18.920 ;
        RECT 85.430 18.840 85.750 19.150 ;
        RECT 87.070 18.840 87.390 19.150 ;
        RECT 87.980 18.840 88.300 19.150 ;
        RECT 89.610 18.920 89.900 19.180 ;
        RECT 89.680 18.700 89.820 18.920 ;
        RECT 91.180 18.840 91.500 19.150 ;
        RECT 92.820 18.840 93.140 19.150 ;
        RECT 93.730 18.840 94.050 19.150 ;
        RECT 1.260 18.560 94.660 18.700 ;
        RECT 1.260 18.500 1.580 18.560 ;
        RECT 2.960 18.100 3.280 18.410 ;
        RECT 3.870 18.100 4.190 18.410 ;
        RECT 7.060 18.320 7.350 18.560 ;
        RECT 5.460 18.010 5.830 18.320 ;
        RECT 8.710 18.100 9.030 18.410 ;
        RECT 9.620 18.100 9.940 18.410 ;
        RECT 12.810 18.320 13.100 18.560 ;
        RECT 11.210 18.010 11.580 18.320 ;
        RECT 14.460 18.100 14.780 18.410 ;
        RECT 15.370 18.100 15.690 18.410 ;
        RECT 18.560 18.320 18.850 18.560 ;
        RECT 16.960 18.010 17.330 18.320 ;
        RECT 20.210 18.100 20.530 18.410 ;
        RECT 21.120 18.100 21.440 18.410 ;
        RECT 24.310 18.320 24.600 18.560 ;
        RECT 22.710 18.010 23.080 18.320 ;
        RECT 25.960 18.100 26.280 18.410 ;
        RECT 26.870 18.100 27.190 18.410 ;
        RECT 30.060 18.320 30.350 18.560 ;
        RECT 28.460 18.010 28.830 18.320 ;
        RECT 31.710 18.100 32.030 18.410 ;
        RECT 32.620 18.100 32.940 18.410 ;
        RECT 35.810 18.320 36.100 18.560 ;
        RECT 34.210 18.010 34.580 18.320 ;
        RECT 37.460 18.100 37.780 18.410 ;
        RECT 38.370 18.100 38.690 18.410 ;
        RECT 41.560 18.320 41.850 18.560 ;
        RECT 39.960 18.010 40.330 18.320 ;
        RECT 43.210 18.100 43.530 18.410 ;
        RECT 44.120 18.100 44.440 18.410 ;
        RECT 47.310 18.320 47.600 18.560 ;
        RECT 45.710 18.010 46.080 18.320 ;
        RECT 48.960 18.100 49.280 18.410 ;
        RECT 49.870 18.100 50.190 18.410 ;
        RECT 53.060 18.320 53.350 18.560 ;
        RECT 51.460 18.010 51.830 18.320 ;
        RECT 54.710 18.100 55.030 18.410 ;
        RECT 55.620 18.100 55.940 18.410 ;
        RECT 58.810 18.320 59.100 18.560 ;
        RECT 57.210 18.010 57.580 18.320 ;
        RECT 60.460 18.100 60.780 18.410 ;
        RECT 61.370 18.100 61.690 18.410 ;
        RECT 64.560 18.320 64.850 18.560 ;
        RECT 62.960 18.010 63.330 18.320 ;
        RECT 66.210 18.100 66.530 18.410 ;
        RECT 67.120 18.100 67.440 18.410 ;
        RECT 70.310 18.320 70.600 18.560 ;
        RECT 68.710 18.010 69.080 18.320 ;
        RECT 71.960 18.100 72.280 18.410 ;
        RECT 72.870 18.100 73.190 18.410 ;
        RECT 76.060 18.320 76.350 18.560 ;
        RECT 74.460 18.010 74.830 18.320 ;
        RECT 77.710 18.100 78.030 18.410 ;
        RECT 78.620 18.100 78.940 18.410 ;
        RECT 81.810 18.320 82.100 18.560 ;
        RECT 80.210 18.010 80.580 18.320 ;
        RECT 83.460 18.100 83.780 18.410 ;
        RECT 84.370 18.100 84.690 18.410 ;
        RECT 87.560 18.320 87.850 18.560 ;
        RECT 85.960 18.010 86.330 18.320 ;
        RECT 89.210 18.100 89.530 18.410 ;
        RECT 90.120 18.100 90.440 18.410 ;
        RECT 93.310 18.320 93.600 18.560 ;
        RECT 91.710 18.010 92.080 18.320 ;
        RECT 3.360 16.510 3.650 16.770 ;
        RECT 1.260 16.290 1.580 16.350 ;
        RECT 3.430 16.290 3.570 16.510 ;
        RECT 4.930 16.430 5.250 16.740 ;
        RECT 6.570 16.430 6.890 16.740 ;
        RECT 7.480 16.430 7.800 16.740 ;
        RECT 9.110 16.510 9.400 16.770 ;
        RECT 9.180 16.290 9.320 16.510 ;
        RECT 10.680 16.430 11.000 16.740 ;
        RECT 12.320 16.430 12.640 16.740 ;
        RECT 13.230 16.430 13.550 16.740 ;
        RECT 14.860 16.510 15.150 16.770 ;
        RECT 14.930 16.290 15.070 16.510 ;
        RECT 16.430 16.430 16.750 16.740 ;
        RECT 18.070 16.430 18.390 16.740 ;
        RECT 18.980 16.430 19.300 16.740 ;
        RECT 20.610 16.510 20.900 16.770 ;
        RECT 20.680 16.290 20.820 16.510 ;
        RECT 22.180 16.430 22.500 16.740 ;
        RECT 23.820 16.430 24.140 16.740 ;
        RECT 24.730 16.430 25.050 16.740 ;
        RECT 26.360 16.510 26.650 16.770 ;
        RECT 26.430 16.290 26.570 16.510 ;
        RECT 27.930 16.430 28.250 16.740 ;
        RECT 29.570 16.430 29.890 16.740 ;
        RECT 30.480 16.430 30.800 16.740 ;
        RECT 32.110 16.510 32.400 16.770 ;
        RECT 32.180 16.290 32.320 16.510 ;
        RECT 33.680 16.430 34.000 16.740 ;
        RECT 35.320 16.430 35.640 16.740 ;
        RECT 36.230 16.430 36.550 16.740 ;
        RECT 37.860 16.510 38.150 16.770 ;
        RECT 37.930 16.290 38.070 16.510 ;
        RECT 39.430 16.430 39.750 16.740 ;
        RECT 41.070 16.430 41.390 16.740 ;
        RECT 41.980 16.430 42.300 16.740 ;
        RECT 43.610 16.510 43.900 16.770 ;
        RECT 43.680 16.290 43.820 16.510 ;
        RECT 45.180 16.430 45.500 16.740 ;
        RECT 46.820 16.430 47.140 16.740 ;
        RECT 47.730 16.430 48.050 16.740 ;
        RECT 49.360 16.510 49.650 16.770 ;
        RECT 49.430 16.290 49.570 16.510 ;
        RECT 50.930 16.430 51.250 16.740 ;
        RECT 52.570 16.430 52.890 16.740 ;
        RECT 53.480 16.430 53.800 16.740 ;
        RECT 55.110 16.510 55.400 16.770 ;
        RECT 55.180 16.290 55.320 16.510 ;
        RECT 56.680 16.430 57.000 16.740 ;
        RECT 58.320 16.430 58.640 16.740 ;
        RECT 59.230 16.430 59.550 16.740 ;
        RECT 60.860 16.510 61.150 16.770 ;
        RECT 60.930 16.290 61.070 16.510 ;
        RECT 62.430 16.430 62.750 16.740 ;
        RECT 64.070 16.430 64.390 16.740 ;
        RECT 64.980 16.430 65.300 16.740 ;
        RECT 66.610 16.510 66.900 16.770 ;
        RECT 66.680 16.290 66.820 16.510 ;
        RECT 68.180 16.430 68.500 16.740 ;
        RECT 69.820 16.430 70.140 16.740 ;
        RECT 70.730 16.430 71.050 16.740 ;
        RECT 72.360 16.510 72.650 16.770 ;
        RECT 72.430 16.290 72.570 16.510 ;
        RECT 73.930 16.430 74.250 16.740 ;
        RECT 75.570 16.430 75.890 16.740 ;
        RECT 76.480 16.430 76.800 16.740 ;
        RECT 78.110 16.510 78.400 16.770 ;
        RECT 78.180 16.290 78.320 16.510 ;
        RECT 79.680 16.430 80.000 16.740 ;
        RECT 81.320 16.430 81.640 16.740 ;
        RECT 82.230 16.430 82.550 16.740 ;
        RECT 83.860 16.510 84.150 16.770 ;
        RECT 83.930 16.290 84.070 16.510 ;
        RECT 85.430 16.430 85.750 16.740 ;
        RECT 87.070 16.430 87.390 16.740 ;
        RECT 87.980 16.430 88.300 16.740 ;
        RECT 89.610 16.510 89.900 16.770 ;
        RECT 89.680 16.290 89.820 16.510 ;
        RECT 91.180 16.430 91.500 16.740 ;
        RECT 92.820 16.430 93.140 16.740 ;
        RECT 93.730 16.430 94.050 16.740 ;
        RECT 1.260 16.150 94.660 16.290 ;
        RECT 1.260 16.090 1.580 16.150 ;
        RECT 2.960 15.690 3.280 16.000 ;
        RECT 3.870 15.690 4.190 16.000 ;
        RECT 7.060 15.910 7.350 16.150 ;
        RECT 5.460 15.600 5.830 15.910 ;
        RECT 8.710 15.690 9.030 16.000 ;
        RECT 9.620 15.690 9.940 16.000 ;
        RECT 12.810 15.910 13.100 16.150 ;
        RECT 11.210 15.600 11.580 15.910 ;
        RECT 14.460 15.690 14.780 16.000 ;
        RECT 15.370 15.690 15.690 16.000 ;
        RECT 18.560 15.910 18.850 16.150 ;
        RECT 16.960 15.600 17.330 15.910 ;
        RECT 20.210 15.690 20.530 16.000 ;
        RECT 21.120 15.690 21.440 16.000 ;
        RECT 24.310 15.910 24.600 16.150 ;
        RECT 22.710 15.600 23.080 15.910 ;
        RECT 25.960 15.690 26.280 16.000 ;
        RECT 26.870 15.690 27.190 16.000 ;
        RECT 30.060 15.910 30.350 16.150 ;
        RECT 28.460 15.600 28.830 15.910 ;
        RECT 31.710 15.690 32.030 16.000 ;
        RECT 32.620 15.690 32.940 16.000 ;
        RECT 35.810 15.910 36.100 16.150 ;
        RECT 34.210 15.600 34.580 15.910 ;
        RECT 37.460 15.690 37.780 16.000 ;
        RECT 38.370 15.690 38.690 16.000 ;
        RECT 41.560 15.910 41.850 16.150 ;
        RECT 39.960 15.600 40.330 15.910 ;
        RECT 43.210 15.690 43.530 16.000 ;
        RECT 44.120 15.690 44.440 16.000 ;
        RECT 47.310 15.910 47.600 16.150 ;
        RECT 45.710 15.600 46.080 15.910 ;
        RECT 48.960 15.690 49.280 16.000 ;
        RECT 49.870 15.690 50.190 16.000 ;
        RECT 53.060 15.910 53.350 16.150 ;
        RECT 51.460 15.600 51.830 15.910 ;
        RECT 54.710 15.690 55.030 16.000 ;
        RECT 55.620 15.690 55.940 16.000 ;
        RECT 58.810 15.910 59.100 16.150 ;
        RECT 57.210 15.600 57.580 15.910 ;
        RECT 60.460 15.690 60.780 16.000 ;
        RECT 61.370 15.690 61.690 16.000 ;
        RECT 64.560 15.910 64.850 16.150 ;
        RECT 62.960 15.600 63.330 15.910 ;
        RECT 66.210 15.690 66.530 16.000 ;
        RECT 67.120 15.690 67.440 16.000 ;
        RECT 70.310 15.910 70.600 16.150 ;
        RECT 68.710 15.600 69.080 15.910 ;
        RECT 71.960 15.690 72.280 16.000 ;
        RECT 72.870 15.690 73.190 16.000 ;
        RECT 76.060 15.910 76.350 16.150 ;
        RECT 74.460 15.600 74.830 15.910 ;
        RECT 77.710 15.690 78.030 16.000 ;
        RECT 78.620 15.690 78.940 16.000 ;
        RECT 81.810 15.910 82.100 16.150 ;
        RECT 80.210 15.600 80.580 15.910 ;
        RECT 83.460 15.690 83.780 16.000 ;
        RECT 84.370 15.690 84.690 16.000 ;
        RECT 87.560 15.910 87.850 16.150 ;
        RECT 85.960 15.600 86.330 15.910 ;
        RECT 89.210 15.690 89.530 16.000 ;
        RECT 90.120 15.690 90.440 16.000 ;
        RECT 93.310 15.910 93.600 16.150 ;
        RECT 91.710 15.600 92.080 15.910 ;
        RECT 3.360 14.100 3.650 14.360 ;
        RECT 1.260 13.880 1.580 13.940 ;
        RECT 3.430 13.880 3.570 14.100 ;
        RECT 4.930 14.020 5.250 14.330 ;
        RECT 6.570 14.020 6.890 14.330 ;
        RECT 7.480 14.020 7.800 14.330 ;
        RECT 9.110 14.100 9.400 14.360 ;
        RECT 9.180 13.880 9.320 14.100 ;
        RECT 10.680 14.020 11.000 14.330 ;
        RECT 12.320 14.020 12.640 14.330 ;
        RECT 13.230 14.020 13.550 14.330 ;
        RECT 14.860 14.100 15.150 14.360 ;
        RECT 14.930 13.880 15.070 14.100 ;
        RECT 16.430 14.020 16.750 14.330 ;
        RECT 18.070 14.020 18.390 14.330 ;
        RECT 18.980 14.020 19.300 14.330 ;
        RECT 20.610 14.100 20.900 14.360 ;
        RECT 20.680 13.880 20.820 14.100 ;
        RECT 22.180 14.020 22.500 14.330 ;
        RECT 23.820 14.020 24.140 14.330 ;
        RECT 24.730 14.020 25.050 14.330 ;
        RECT 26.360 14.100 26.650 14.360 ;
        RECT 26.430 13.880 26.570 14.100 ;
        RECT 27.930 14.020 28.250 14.330 ;
        RECT 29.570 14.020 29.890 14.330 ;
        RECT 30.480 14.020 30.800 14.330 ;
        RECT 32.110 14.100 32.400 14.360 ;
        RECT 32.180 13.880 32.320 14.100 ;
        RECT 33.680 14.020 34.000 14.330 ;
        RECT 35.320 14.020 35.640 14.330 ;
        RECT 36.230 14.020 36.550 14.330 ;
        RECT 37.860 14.100 38.150 14.360 ;
        RECT 37.930 13.880 38.070 14.100 ;
        RECT 39.430 14.020 39.750 14.330 ;
        RECT 41.070 14.020 41.390 14.330 ;
        RECT 41.980 14.020 42.300 14.330 ;
        RECT 43.610 14.100 43.900 14.360 ;
        RECT 43.680 13.880 43.820 14.100 ;
        RECT 45.180 14.020 45.500 14.330 ;
        RECT 46.820 14.020 47.140 14.330 ;
        RECT 47.730 14.020 48.050 14.330 ;
        RECT 49.360 14.100 49.650 14.360 ;
        RECT 49.430 13.880 49.570 14.100 ;
        RECT 50.930 14.020 51.250 14.330 ;
        RECT 52.570 14.020 52.890 14.330 ;
        RECT 53.480 14.020 53.800 14.330 ;
        RECT 55.110 14.100 55.400 14.360 ;
        RECT 55.180 13.880 55.320 14.100 ;
        RECT 56.680 14.020 57.000 14.330 ;
        RECT 58.320 14.020 58.640 14.330 ;
        RECT 59.230 14.020 59.550 14.330 ;
        RECT 60.860 14.100 61.150 14.360 ;
        RECT 60.930 13.880 61.070 14.100 ;
        RECT 62.430 14.020 62.750 14.330 ;
        RECT 64.070 14.020 64.390 14.330 ;
        RECT 64.980 14.020 65.300 14.330 ;
        RECT 66.610 14.100 66.900 14.360 ;
        RECT 66.680 13.880 66.820 14.100 ;
        RECT 68.180 14.020 68.500 14.330 ;
        RECT 69.820 14.020 70.140 14.330 ;
        RECT 70.730 14.020 71.050 14.330 ;
        RECT 72.360 14.100 72.650 14.360 ;
        RECT 72.430 13.880 72.570 14.100 ;
        RECT 73.930 14.020 74.250 14.330 ;
        RECT 75.570 14.020 75.890 14.330 ;
        RECT 76.480 14.020 76.800 14.330 ;
        RECT 78.110 14.100 78.400 14.360 ;
        RECT 78.180 13.880 78.320 14.100 ;
        RECT 79.680 14.020 80.000 14.330 ;
        RECT 81.320 14.020 81.640 14.330 ;
        RECT 82.230 14.020 82.550 14.330 ;
        RECT 83.860 14.100 84.150 14.360 ;
        RECT 83.930 13.880 84.070 14.100 ;
        RECT 85.430 14.020 85.750 14.330 ;
        RECT 87.070 14.020 87.390 14.330 ;
        RECT 87.980 14.020 88.300 14.330 ;
        RECT 89.610 14.100 89.900 14.360 ;
        RECT 89.680 13.880 89.820 14.100 ;
        RECT 91.180 14.020 91.500 14.330 ;
        RECT 92.820 14.020 93.140 14.330 ;
        RECT 93.730 14.020 94.050 14.330 ;
        RECT 1.260 13.740 94.660 13.880 ;
        RECT 1.260 13.680 1.580 13.740 ;
        RECT 2.960 13.280 3.280 13.590 ;
        RECT 3.870 13.280 4.190 13.590 ;
        RECT 7.060 13.500 7.350 13.740 ;
        RECT 5.460 13.190 5.830 13.500 ;
        RECT 8.710 13.280 9.030 13.590 ;
        RECT 9.620 13.280 9.940 13.590 ;
        RECT 12.810 13.500 13.100 13.740 ;
        RECT 11.210 13.190 11.580 13.500 ;
        RECT 14.460 13.280 14.780 13.590 ;
        RECT 15.370 13.280 15.690 13.590 ;
        RECT 18.560 13.500 18.850 13.740 ;
        RECT 16.960 13.190 17.330 13.500 ;
        RECT 20.210 13.280 20.530 13.590 ;
        RECT 21.120 13.280 21.440 13.590 ;
        RECT 24.310 13.500 24.600 13.740 ;
        RECT 22.710 13.190 23.080 13.500 ;
        RECT 25.960 13.280 26.280 13.590 ;
        RECT 26.870 13.280 27.190 13.590 ;
        RECT 30.060 13.500 30.350 13.740 ;
        RECT 28.460 13.190 28.830 13.500 ;
        RECT 31.710 13.280 32.030 13.590 ;
        RECT 32.620 13.280 32.940 13.590 ;
        RECT 35.810 13.500 36.100 13.740 ;
        RECT 34.210 13.190 34.580 13.500 ;
        RECT 37.460 13.280 37.780 13.590 ;
        RECT 38.370 13.280 38.690 13.590 ;
        RECT 41.560 13.500 41.850 13.740 ;
        RECT 39.960 13.190 40.330 13.500 ;
        RECT 43.210 13.280 43.530 13.590 ;
        RECT 44.120 13.280 44.440 13.590 ;
        RECT 47.310 13.500 47.600 13.740 ;
        RECT 45.710 13.190 46.080 13.500 ;
        RECT 48.960 13.280 49.280 13.590 ;
        RECT 49.870 13.280 50.190 13.590 ;
        RECT 53.060 13.500 53.350 13.740 ;
        RECT 51.460 13.190 51.830 13.500 ;
        RECT 54.710 13.280 55.030 13.590 ;
        RECT 55.620 13.280 55.940 13.590 ;
        RECT 58.810 13.500 59.100 13.740 ;
        RECT 57.210 13.190 57.580 13.500 ;
        RECT 60.460 13.280 60.780 13.590 ;
        RECT 61.370 13.280 61.690 13.590 ;
        RECT 64.560 13.500 64.850 13.740 ;
        RECT 62.960 13.190 63.330 13.500 ;
        RECT 66.210 13.280 66.530 13.590 ;
        RECT 67.120 13.280 67.440 13.590 ;
        RECT 70.310 13.500 70.600 13.740 ;
        RECT 68.710 13.190 69.080 13.500 ;
        RECT 71.960 13.280 72.280 13.590 ;
        RECT 72.870 13.280 73.190 13.590 ;
        RECT 76.060 13.500 76.350 13.740 ;
        RECT 74.460 13.190 74.830 13.500 ;
        RECT 77.710 13.280 78.030 13.590 ;
        RECT 78.620 13.280 78.940 13.590 ;
        RECT 81.810 13.500 82.100 13.740 ;
        RECT 80.210 13.190 80.580 13.500 ;
        RECT 83.460 13.280 83.780 13.590 ;
        RECT 84.370 13.280 84.690 13.590 ;
        RECT 87.560 13.500 87.850 13.740 ;
        RECT 85.960 13.190 86.330 13.500 ;
        RECT 89.210 13.280 89.530 13.590 ;
        RECT 90.120 13.280 90.440 13.590 ;
        RECT 93.310 13.500 93.600 13.740 ;
        RECT 91.710 13.190 92.080 13.500 ;
        RECT 3.360 11.690 3.650 11.950 ;
        RECT 1.250 11.470 1.570 11.530 ;
        RECT 3.430 11.470 3.570 11.690 ;
        RECT 4.930 11.610 5.250 11.920 ;
        RECT 6.570 11.610 6.890 11.920 ;
        RECT 7.480 11.610 7.800 11.920 ;
        RECT 9.110 11.690 9.400 11.950 ;
        RECT 9.180 11.470 9.320 11.690 ;
        RECT 10.680 11.610 11.000 11.920 ;
        RECT 12.320 11.610 12.640 11.920 ;
        RECT 13.230 11.610 13.550 11.920 ;
        RECT 14.860 11.690 15.150 11.950 ;
        RECT 14.930 11.470 15.070 11.690 ;
        RECT 16.430 11.610 16.750 11.920 ;
        RECT 18.070 11.610 18.390 11.920 ;
        RECT 18.980 11.610 19.300 11.920 ;
        RECT 20.610 11.690 20.900 11.950 ;
        RECT 20.680 11.470 20.820 11.690 ;
        RECT 22.180 11.610 22.500 11.920 ;
        RECT 23.820 11.610 24.140 11.920 ;
        RECT 24.730 11.610 25.050 11.920 ;
        RECT 26.360 11.690 26.650 11.950 ;
        RECT 26.430 11.470 26.570 11.690 ;
        RECT 27.930 11.610 28.250 11.920 ;
        RECT 29.570 11.610 29.890 11.920 ;
        RECT 30.480 11.610 30.800 11.920 ;
        RECT 32.110 11.690 32.400 11.950 ;
        RECT 32.180 11.470 32.320 11.690 ;
        RECT 33.680 11.610 34.000 11.920 ;
        RECT 35.320 11.610 35.640 11.920 ;
        RECT 36.230 11.610 36.550 11.920 ;
        RECT 37.860 11.690 38.150 11.950 ;
        RECT 37.930 11.470 38.070 11.690 ;
        RECT 39.430 11.610 39.750 11.920 ;
        RECT 41.070 11.610 41.390 11.920 ;
        RECT 41.980 11.610 42.300 11.920 ;
        RECT 43.610 11.690 43.900 11.950 ;
        RECT 43.680 11.470 43.820 11.690 ;
        RECT 45.180 11.610 45.500 11.920 ;
        RECT 46.820 11.610 47.140 11.920 ;
        RECT 47.730 11.610 48.050 11.920 ;
        RECT 49.360 11.690 49.650 11.950 ;
        RECT 49.430 11.470 49.570 11.690 ;
        RECT 50.930 11.610 51.250 11.920 ;
        RECT 52.570 11.610 52.890 11.920 ;
        RECT 53.480 11.610 53.800 11.920 ;
        RECT 55.110 11.690 55.400 11.950 ;
        RECT 55.180 11.470 55.320 11.690 ;
        RECT 56.680 11.610 57.000 11.920 ;
        RECT 58.320 11.610 58.640 11.920 ;
        RECT 59.230 11.610 59.550 11.920 ;
        RECT 60.860 11.690 61.150 11.950 ;
        RECT 60.930 11.470 61.070 11.690 ;
        RECT 62.430 11.610 62.750 11.920 ;
        RECT 64.070 11.610 64.390 11.920 ;
        RECT 64.980 11.610 65.300 11.920 ;
        RECT 66.610 11.690 66.900 11.950 ;
        RECT 66.680 11.470 66.820 11.690 ;
        RECT 68.180 11.610 68.500 11.920 ;
        RECT 69.820 11.610 70.140 11.920 ;
        RECT 70.730 11.610 71.050 11.920 ;
        RECT 72.360 11.690 72.650 11.950 ;
        RECT 72.430 11.470 72.570 11.690 ;
        RECT 73.930 11.610 74.250 11.920 ;
        RECT 75.570 11.610 75.890 11.920 ;
        RECT 76.480 11.610 76.800 11.920 ;
        RECT 78.110 11.690 78.400 11.950 ;
        RECT 78.180 11.470 78.320 11.690 ;
        RECT 79.680 11.610 80.000 11.920 ;
        RECT 81.320 11.610 81.640 11.920 ;
        RECT 82.230 11.610 82.550 11.920 ;
        RECT 83.860 11.690 84.150 11.950 ;
        RECT 83.930 11.470 84.070 11.690 ;
        RECT 85.430 11.610 85.750 11.920 ;
        RECT 87.070 11.610 87.390 11.920 ;
        RECT 87.980 11.610 88.300 11.920 ;
        RECT 89.610 11.690 89.900 11.950 ;
        RECT 89.680 11.470 89.820 11.690 ;
        RECT 91.180 11.610 91.500 11.920 ;
        RECT 92.820 11.610 93.140 11.920 ;
        RECT 93.730 11.610 94.050 11.920 ;
        RECT 1.250 11.330 94.660 11.470 ;
        RECT 1.250 11.270 1.570 11.330 ;
        RECT 2.960 10.870 3.280 11.180 ;
        RECT 3.870 10.870 4.190 11.180 ;
        RECT 7.060 11.090 7.350 11.330 ;
        RECT 5.460 10.780 5.830 11.090 ;
        RECT 8.710 10.870 9.030 11.180 ;
        RECT 9.620 10.870 9.940 11.180 ;
        RECT 12.810 11.090 13.100 11.330 ;
        RECT 11.210 10.780 11.580 11.090 ;
        RECT 14.460 10.870 14.780 11.180 ;
        RECT 15.370 10.870 15.690 11.180 ;
        RECT 18.560 11.090 18.850 11.330 ;
        RECT 16.960 10.780 17.330 11.090 ;
        RECT 20.210 10.870 20.530 11.180 ;
        RECT 21.120 10.870 21.440 11.180 ;
        RECT 24.310 11.090 24.600 11.330 ;
        RECT 22.710 10.780 23.080 11.090 ;
        RECT 25.960 10.870 26.280 11.180 ;
        RECT 26.870 10.870 27.190 11.180 ;
        RECT 30.060 11.090 30.350 11.330 ;
        RECT 28.460 10.780 28.830 11.090 ;
        RECT 31.710 10.870 32.030 11.180 ;
        RECT 32.620 10.870 32.940 11.180 ;
        RECT 35.810 11.090 36.100 11.330 ;
        RECT 34.210 10.780 34.580 11.090 ;
        RECT 37.460 10.870 37.780 11.180 ;
        RECT 38.370 10.870 38.690 11.180 ;
        RECT 41.560 11.090 41.850 11.330 ;
        RECT 39.960 10.780 40.330 11.090 ;
        RECT 43.210 10.870 43.530 11.180 ;
        RECT 44.120 10.870 44.440 11.180 ;
        RECT 47.310 11.090 47.600 11.330 ;
        RECT 45.710 10.780 46.080 11.090 ;
        RECT 48.960 10.870 49.280 11.180 ;
        RECT 49.870 10.870 50.190 11.180 ;
        RECT 53.060 11.090 53.350 11.330 ;
        RECT 51.460 10.780 51.830 11.090 ;
        RECT 54.710 10.870 55.030 11.180 ;
        RECT 55.620 10.870 55.940 11.180 ;
        RECT 58.810 11.090 59.100 11.330 ;
        RECT 57.210 10.780 57.580 11.090 ;
        RECT 60.460 10.870 60.780 11.180 ;
        RECT 61.370 10.870 61.690 11.180 ;
        RECT 64.560 11.090 64.850 11.330 ;
        RECT 62.960 10.780 63.330 11.090 ;
        RECT 66.210 10.870 66.530 11.180 ;
        RECT 67.120 10.870 67.440 11.180 ;
        RECT 70.310 11.090 70.600 11.330 ;
        RECT 68.710 10.780 69.080 11.090 ;
        RECT 71.960 10.870 72.280 11.180 ;
        RECT 72.870 10.870 73.190 11.180 ;
        RECT 76.060 11.090 76.350 11.330 ;
        RECT 74.460 10.780 74.830 11.090 ;
        RECT 77.710 10.870 78.030 11.180 ;
        RECT 78.620 10.870 78.940 11.180 ;
        RECT 81.810 11.090 82.100 11.330 ;
        RECT 80.210 10.780 80.580 11.090 ;
        RECT 83.460 10.870 83.780 11.180 ;
        RECT 84.370 10.870 84.690 11.180 ;
        RECT 87.560 11.090 87.850 11.330 ;
        RECT 85.960 10.780 86.330 11.090 ;
        RECT 89.210 10.870 89.530 11.180 ;
        RECT 90.120 10.870 90.440 11.180 ;
        RECT 93.310 11.090 93.600 11.330 ;
        RECT 91.710 10.780 92.080 11.090 ;
        RECT 3.360 9.280 3.650 9.540 ;
        RECT 1.260 9.060 1.580 9.120 ;
        RECT 3.430 9.060 3.570 9.280 ;
        RECT 4.930 9.200 5.250 9.510 ;
        RECT 6.570 9.200 6.890 9.510 ;
        RECT 7.480 9.200 7.800 9.510 ;
        RECT 9.110 9.280 9.400 9.540 ;
        RECT 9.180 9.060 9.320 9.280 ;
        RECT 10.680 9.200 11.000 9.510 ;
        RECT 12.320 9.200 12.640 9.510 ;
        RECT 13.230 9.200 13.550 9.510 ;
        RECT 14.860 9.280 15.150 9.540 ;
        RECT 14.930 9.060 15.070 9.280 ;
        RECT 16.430 9.200 16.750 9.510 ;
        RECT 18.070 9.200 18.390 9.510 ;
        RECT 18.980 9.200 19.300 9.510 ;
        RECT 20.610 9.280 20.900 9.540 ;
        RECT 20.680 9.060 20.820 9.280 ;
        RECT 22.180 9.200 22.500 9.510 ;
        RECT 23.820 9.200 24.140 9.510 ;
        RECT 24.730 9.200 25.050 9.510 ;
        RECT 26.360 9.280 26.650 9.540 ;
        RECT 26.430 9.060 26.570 9.280 ;
        RECT 27.930 9.200 28.250 9.510 ;
        RECT 29.570 9.200 29.890 9.510 ;
        RECT 30.480 9.200 30.800 9.510 ;
        RECT 32.110 9.280 32.400 9.540 ;
        RECT 32.180 9.060 32.320 9.280 ;
        RECT 33.680 9.200 34.000 9.510 ;
        RECT 35.320 9.200 35.640 9.510 ;
        RECT 36.230 9.200 36.550 9.510 ;
        RECT 37.860 9.280 38.150 9.540 ;
        RECT 37.930 9.060 38.070 9.280 ;
        RECT 39.430 9.200 39.750 9.510 ;
        RECT 41.070 9.200 41.390 9.510 ;
        RECT 41.980 9.200 42.300 9.510 ;
        RECT 43.610 9.280 43.900 9.540 ;
        RECT 43.680 9.060 43.820 9.280 ;
        RECT 45.180 9.200 45.500 9.510 ;
        RECT 46.820 9.200 47.140 9.510 ;
        RECT 47.730 9.200 48.050 9.510 ;
        RECT 49.360 9.280 49.650 9.540 ;
        RECT 49.430 9.060 49.570 9.280 ;
        RECT 50.930 9.200 51.250 9.510 ;
        RECT 52.570 9.200 52.890 9.510 ;
        RECT 53.480 9.200 53.800 9.510 ;
        RECT 55.110 9.280 55.400 9.540 ;
        RECT 55.180 9.060 55.320 9.280 ;
        RECT 56.680 9.200 57.000 9.510 ;
        RECT 58.320 9.200 58.640 9.510 ;
        RECT 59.230 9.200 59.550 9.510 ;
        RECT 60.860 9.280 61.150 9.540 ;
        RECT 60.930 9.060 61.070 9.280 ;
        RECT 62.430 9.200 62.750 9.510 ;
        RECT 64.070 9.200 64.390 9.510 ;
        RECT 64.980 9.200 65.300 9.510 ;
        RECT 66.610 9.280 66.900 9.540 ;
        RECT 66.680 9.060 66.820 9.280 ;
        RECT 68.180 9.200 68.500 9.510 ;
        RECT 69.820 9.200 70.140 9.510 ;
        RECT 70.730 9.200 71.050 9.510 ;
        RECT 72.360 9.280 72.650 9.540 ;
        RECT 72.430 9.060 72.570 9.280 ;
        RECT 73.930 9.200 74.250 9.510 ;
        RECT 75.570 9.200 75.890 9.510 ;
        RECT 76.480 9.200 76.800 9.510 ;
        RECT 78.110 9.280 78.400 9.540 ;
        RECT 78.180 9.060 78.320 9.280 ;
        RECT 79.680 9.200 80.000 9.510 ;
        RECT 81.320 9.200 81.640 9.510 ;
        RECT 82.230 9.200 82.550 9.510 ;
        RECT 83.860 9.280 84.150 9.540 ;
        RECT 83.930 9.060 84.070 9.280 ;
        RECT 85.430 9.200 85.750 9.510 ;
        RECT 87.070 9.200 87.390 9.510 ;
        RECT 87.980 9.200 88.300 9.510 ;
        RECT 89.610 9.280 89.900 9.540 ;
        RECT 89.680 9.060 89.820 9.280 ;
        RECT 91.180 9.200 91.500 9.510 ;
        RECT 92.820 9.200 93.140 9.510 ;
        RECT 93.730 9.200 94.050 9.510 ;
        RECT 1.260 8.920 94.660 9.060 ;
        RECT 1.260 8.860 1.580 8.920 ;
        RECT 7.140 8.630 7.280 8.920 ;
        RECT 12.890 8.630 13.030 8.920 ;
        RECT 18.640 8.630 18.780 8.920 ;
        RECT 24.390 8.630 24.530 8.920 ;
        RECT 30.140 8.630 30.280 8.920 ;
        RECT 35.890 8.630 36.030 8.920 ;
        RECT 41.640 8.630 41.780 8.920 ;
        RECT 47.390 8.630 47.530 8.920 ;
        RECT 53.140 8.630 53.280 8.920 ;
        RECT 58.890 8.630 59.030 8.920 ;
        RECT 64.640 8.630 64.780 8.920 ;
        RECT 70.390 8.630 70.530 8.920 ;
        RECT 76.140 8.630 76.280 8.920 ;
        RECT 81.890 8.630 82.030 8.920 ;
        RECT 87.640 8.630 87.780 8.920 ;
        RECT 93.390 8.630 93.530 8.920 ;
        RECT 7.060 8.380 7.350 8.630 ;
        RECT 12.810 8.380 13.100 8.630 ;
        RECT 18.560 8.380 18.850 8.630 ;
        RECT 24.310 8.380 24.600 8.630 ;
        RECT 30.060 8.380 30.350 8.630 ;
        RECT 35.810 8.380 36.100 8.630 ;
        RECT 41.560 8.380 41.850 8.630 ;
        RECT 47.310 8.380 47.600 8.630 ;
        RECT 53.060 8.380 53.350 8.630 ;
        RECT 58.810 8.380 59.100 8.630 ;
        RECT 64.560 8.380 64.850 8.630 ;
        RECT 70.310 8.380 70.600 8.630 ;
        RECT 76.060 8.380 76.350 8.630 ;
        RECT 81.810 8.380 82.100 8.630 ;
        RECT 87.560 8.380 87.850 8.630 ;
        RECT 93.310 8.380 93.600 8.630 ;
        RECT 2.960 8.050 3.280 8.360 ;
        RECT 3.870 8.050 4.190 8.360 ;
        RECT 5.460 7.960 5.830 8.270 ;
        RECT 8.710 8.050 9.030 8.360 ;
        RECT 9.620 8.050 9.940 8.360 ;
        RECT 11.210 7.960 11.580 8.270 ;
        RECT 14.460 8.050 14.780 8.360 ;
        RECT 15.370 8.050 15.690 8.360 ;
        RECT 16.960 7.960 17.330 8.270 ;
        RECT 20.210 8.050 20.530 8.360 ;
        RECT 21.120 8.050 21.440 8.360 ;
        RECT 22.710 7.960 23.080 8.270 ;
        RECT 25.960 8.050 26.280 8.360 ;
        RECT 26.870 8.050 27.190 8.360 ;
        RECT 28.460 7.960 28.830 8.270 ;
        RECT 31.710 8.050 32.030 8.360 ;
        RECT 32.620 8.050 32.940 8.360 ;
        RECT 34.210 7.960 34.580 8.270 ;
        RECT 37.460 8.050 37.780 8.360 ;
        RECT 38.370 8.050 38.690 8.360 ;
        RECT 39.960 7.960 40.330 8.270 ;
        RECT 43.210 8.050 43.530 8.360 ;
        RECT 44.120 8.050 44.440 8.360 ;
        RECT 45.710 7.960 46.080 8.270 ;
        RECT 48.960 8.050 49.280 8.360 ;
        RECT 49.870 8.050 50.190 8.360 ;
        RECT 51.460 7.960 51.830 8.270 ;
        RECT 54.710 8.050 55.030 8.360 ;
        RECT 55.620 8.050 55.940 8.360 ;
        RECT 57.210 7.960 57.580 8.270 ;
        RECT 60.460 8.050 60.780 8.360 ;
        RECT 61.370 8.050 61.690 8.360 ;
        RECT 62.960 7.960 63.330 8.270 ;
        RECT 66.210 8.050 66.530 8.360 ;
        RECT 67.120 8.050 67.440 8.360 ;
        RECT 68.710 7.960 69.080 8.270 ;
        RECT 71.960 8.050 72.280 8.360 ;
        RECT 72.870 8.050 73.190 8.360 ;
        RECT 74.460 7.960 74.830 8.270 ;
        RECT 77.710 8.050 78.030 8.360 ;
        RECT 78.620 8.050 78.940 8.360 ;
        RECT 80.210 7.960 80.580 8.270 ;
        RECT 83.460 8.050 83.780 8.360 ;
        RECT 84.370 8.050 84.690 8.360 ;
        RECT 85.960 7.960 86.330 8.270 ;
        RECT 89.210 8.050 89.530 8.360 ;
        RECT 90.120 8.050 90.440 8.360 ;
        RECT 91.710 7.960 92.080 8.270 ;
        RECT 3.360 6.460 3.650 6.720 ;
        RECT 1.250 6.240 1.570 6.300 ;
        RECT 3.430 6.240 3.570 6.460 ;
        RECT 4.930 6.380 5.250 6.690 ;
        RECT 6.570 6.380 6.890 6.690 ;
        RECT 7.480 6.380 7.800 6.690 ;
        RECT 9.110 6.460 9.400 6.720 ;
        RECT 9.180 6.240 9.320 6.460 ;
        RECT 10.680 6.380 11.000 6.690 ;
        RECT 12.320 6.380 12.640 6.690 ;
        RECT 13.230 6.380 13.550 6.690 ;
        RECT 14.860 6.460 15.150 6.720 ;
        RECT 14.930 6.240 15.070 6.460 ;
        RECT 16.430 6.380 16.750 6.690 ;
        RECT 18.070 6.380 18.390 6.690 ;
        RECT 18.980 6.380 19.300 6.690 ;
        RECT 20.610 6.460 20.900 6.720 ;
        RECT 20.680 6.240 20.820 6.460 ;
        RECT 22.180 6.380 22.500 6.690 ;
        RECT 23.820 6.380 24.140 6.690 ;
        RECT 24.730 6.380 25.050 6.690 ;
        RECT 26.360 6.460 26.650 6.720 ;
        RECT 26.430 6.240 26.570 6.460 ;
        RECT 27.930 6.380 28.250 6.690 ;
        RECT 29.570 6.380 29.890 6.690 ;
        RECT 30.480 6.380 30.800 6.690 ;
        RECT 32.110 6.460 32.400 6.720 ;
        RECT 32.180 6.240 32.320 6.460 ;
        RECT 33.680 6.380 34.000 6.690 ;
        RECT 35.320 6.380 35.640 6.690 ;
        RECT 36.230 6.380 36.550 6.690 ;
        RECT 37.860 6.460 38.150 6.720 ;
        RECT 37.930 6.240 38.070 6.460 ;
        RECT 39.430 6.380 39.750 6.690 ;
        RECT 41.070 6.380 41.390 6.690 ;
        RECT 41.980 6.380 42.300 6.690 ;
        RECT 43.610 6.460 43.900 6.720 ;
        RECT 43.680 6.240 43.820 6.460 ;
        RECT 45.180 6.380 45.500 6.690 ;
        RECT 46.820 6.380 47.140 6.690 ;
        RECT 47.730 6.380 48.050 6.690 ;
        RECT 49.360 6.460 49.650 6.720 ;
        RECT 49.430 6.240 49.570 6.460 ;
        RECT 50.930 6.380 51.250 6.690 ;
        RECT 52.570 6.380 52.890 6.690 ;
        RECT 53.480 6.380 53.800 6.690 ;
        RECT 55.110 6.460 55.400 6.720 ;
        RECT 55.180 6.240 55.320 6.460 ;
        RECT 56.680 6.380 57.000 6.690 ;
        RECT 58.320 6.380 58.640 6.690 ;
        RECT 59.230 6.380 59.550 6.690 ;
        RECT 60.860 6.460 61.150 6.720 ;
        RECT 60.930 6.240 61.070 6.460 ;
        RECT 62.430 6.380 62.750 6.690 ;
        RECT 64.070 6.380 64.390 6.690 ;
        RECT 64.980 6.380 65.300 6.690 ;
        RECT 66.610 6.460 66.900 6.720 ;
        RECT 66.680 6.240 66.820 6.460 ;
        RECT 68.180 6.380 68.500 6.690 ;
        RECT 69.820 6.380 70.140 6.690 ;
        RECT 70.730 6.380 71.050 6.690 ;
        RECT 72.360 6.460 72.650 6.720 ;
        RECT 72.430 6.240 72.570 6.460 ;
        RECT 73.930 6.380 74.250 6.690 ;
        RECT 75.570 6.380 75.890 6.690 ;
        RECT 76.480 6.380 76.800 6.690 ;
        RECT 78.110 6.460 78.400 6.720 ;
        RECT 78.180 6.240 78.320 6.460 ;
        RECT 79.680 6.380 80.000 6.690 ;
        RECT 81.320 6.380 81.640 6.690 ;
        RECT 82.230 6.380 82.550 6.690 ;
        RECT 83.860 6.460 84.150 6.720 ;
        RECT 83.930 6.240 84.070 6.460 ;
        RECT 85.430 6.380 85.750 6.690 ;
        RECT 87.070 6.380 87.390 6.690 ;
        RECT 87.980 6.380 88.300 6.690 ;
        RECT 89.610 6.460 89.900 6.720 ;
        RECT 89.680 6.240 89.820 6.460 ;
        RECT 91.180 6.380 91.500 6.690 ;
        RECT 92.820 6.380 93.140 6.690 ;
        RECT 93.730 6.380 94.050 6.690 ;
        RECT 1.250 6.100 94.660 6.240 ;
        RECT 1.250 6.040 1.570 6.100 ;
        RECT 2.960 5.640 3.280 5.950 ;
        RECT 3.870 5.640 4.190 5.950 ;
        RECT 7.060 5.860 7.350 6.100 ;
        RECT 5.460 5.550 5.830 5.860 ;
        RECT 8.710 5.640 9.030 5.950 ;
        RECT 9.620 5.640 9.940 5.950 ;
        RECT 12.810 5.860 13.100 6.100 ;
        RECT 11.210 5.550 11.580 5.860 ;
        RECT 14.460 5.640 14.780 5.950 ;
        RECT 15.370 5.640 15.690 5.950 ;
        RECT 18.560 5.860 18.850 6.100 ;
        RECT 16.960 5.550 17.330 5.860 ;
        RECT 20.210 5.640 20.530 5.950 ;
        RECT 21.120 5.640 21.440 5.950 ;
        RECT 24.310 5.860 24.600 6.100 ;
        RECT 22.710 5.550 23.080 5.860 ;
        RECT 25.960 5.640 26.280 5.950 ;
        RECT 26.870 5.640 27.190 5.950 ;
        RECT 30.060 5.860 30.350 6.100 ;
        RECT 28.460 5.550 28.830 5.860 ;
        RECT 31.710 5.640 32.030 5.950 ;
        RECT 32.620 5.640 32.940 5.950 ;
        RECT 35.810 5.860 36.100 6.100 ;
        RECT 34.210 5.550 34.580 5.860 ;
        RECT 37.460 5.640 37.780 5.950 ;
        RECT 38.370 5.640 38.690 5.950 ;
        RECT 41.560 5.860 41.850 6.100 ;
        RECT 39.960 5.550 40.330 5.860 ;
        RECT 43.210 5.640 43.530 5.950 ;
        RECT 44.120 5.640 44.440 5.950 ;
        RECT 47.310 5.860 47.600 6.100 ;
        RECT 45.710 5.550 46.080 5.860 ;
        RECT 48.960 5.640 49.280 5.950 ;
        RECT 49.870 5.640 50.190 5.950 ;
        RECT 53.060 5.860 53.350 6.100 ;
        RECT 51.460 5.550 51.830 5.860 ;
        RECT 54.710 5.640 55.030 5.950 ;
        RECT 55.620 5.640 55.940 5.950 ;
        RECT 58.810 5.860 59.100 6.100 ;
        RECT 57.210 5.550 57.580 5.860 ;
        RECT 60.460 5.640 60.780 5.950 ;
        RECT 61.370 5.640 61.690 5.950 ;
        RECT 64.560 5.860 64.850 6.100 ;
        RECT 62.960 5.550 63.330 5.860 ;
        RECT 66.210 5.640 66.530 5.950 ;
        RECT 67.120 5.640 67.440 5.950 ;
        RECT 70.310 5.860 70.600 6.100 ;
        RECT 68.710 5.550 69.080 5.860 ;
        RECT 71.960 5.640 72.280 5.950 ;
        RECT 72.870 5.640 73.190 5.950 ;
        RECT 76.060 5.860 76.350 6.100 ;
        RECT 74.460 5.550 74.830 5.860 ;
        RECT 77.710 5.640 78.030 5.950 ;
        RECT 78.620 5.640 78.940 5.950 ;
        RECT 81.810 5.860 82.100 6.100 ;
        RECT 80.210 5.550 80.580 5.860 ;
        RECT 83.460 5.640 83.780 5.950 ;
        RECT 84.370 5.640 84.690 5.950 ;
        RECT 87.560 5.860 87.850 6.100 ;
        RECT 85.960 5.550 86.330 5.860 ;
        RECT 89.210 5.640 89.530 5.950 ;
        RECT 90.120 5.640 90.440 5.950 ;
        RECT 93.310 5.860 93.600 6.100 ;
        RECT 91.710 5.550 92.080 5.860 ;
        RECT 3.360 4.050 3.650 4.310 ;
        RECT 1.270 3.830 1.590 3.890 ;
        RECT 3.430 3.830 3.570 4.050 ;
        RECT 4.930 3.970 5.250 4.280 ;
        RECT 6.570 3.970 6.890 4.280 ;
        RECT 7.480 3.970 7.800 4.280 ;
        RECT 9.110 4.050 9.400 4.310 ;
        RECT 9.180 3.830 9.320 4.050 ;
        RECT 10.680 3.970 11.000 4.280 ;
        RECT 12.320 3.970 12.640 4.280 ;
        RECT 13.230 3.970 13.550 4.280 ;
        RECT 14.860 4.050 15.150 4.310 ;
        RECT 14.930 3.830 15.070 4.050 ;
        RECT 16.430 3.970 16.750 4.280 ;
        RECT 18.070 3.970 18.390 4.280 ;
        RECT 18.980 3.970 19.300 4.280 ;
        RECT 20.610 4.050 20.900 4.310 ;
        RECT 20.680 3.830 20.820 4.050 ;
        RECT 22.180 3.970 22.500 4.280 ;
        RECT 23.820 3.970 24.140 4.280 ;
        RECT 24.730 3.970 25.050 4.280 ;
        RECT 26.360 4.050 26.650 4.310 ;
        RECT 26.430 3.830 26.570 4.050 ;
        RECT 27.930 3.970 28.250 4.280 ;
        RECT 29.570 3.970 29.890 4.280 ;
        RECT 30.480 3.970 30.800 4.280 ;
        RECT 32.110 4.050 32.400 4.310 ;
        RECT 32.180 3.830 32.320 4.050 ;
        RECT 33.680 3.970 34.000 4.280 ;
        RECT 35.320 3.970 35.640 4.280 ;
        RECT 36.230 3.970 36.550 4.280 ;
        RECT 37.860 4.050 38.150 4.310 ;
        RECT 37.930 3.830 38.070 4.050 ;
        RECT 39.430 3.970 39.750 4.280 ;
        RECT 41.070 3.970 41.390 4.280 ;
        RECT 41.980 3.970 42.300 4.280 ;
        RECT 43.610 4.050 43.900 4.310 ;
        RECT 43.680 3.830 43.820 4.050 ;
        RECT 45.180 3.970 45.500 4.280 ;
        RECT 46.820 3.970 47.140 4.280 ;
        RECT 47.730 3.970 48.050 4.280 ;
        RECT 49.360 4.050 49.650 4.310 ;
        RECT 49.430 3.830 49.570 4.050 ;
        RECT 50.930 3.970 51.250 4.280 ;
        RECT 52.570 3.970 52.890 4.280 ;
        RECT 53.480 3.970 53.800 4.280 ;
        RECT 55.110 4.050 55.400 4.310 ;
        RECT 55.180 3.830 55.320 4.050 ;
        RECT 56.680 3.970 57.000 4.280 ;
        RECT 58.320 3.970 58.640 4.280 ;
        RECT 59.230 3.970 59.550 4.280 ;
        RECT 60.860 4.050 61.150 4.310 ;
        RECT 60.930 3.830 61.070 4.050 ;
        RECT 62.430 3.970 62.750 4.280 ;
        RECT 64.070 3.970 64.390 4.280 ;
        RECT 64.980 3.970 65.300 4.280 ;
        RECT 66.610 4.050 66.900 4.310 ;
        RECT 66.680 3.830 66.820 4.050 ;
        RECT 68.180 3.970 68.500 4.280 ;
        RECT 69.820 3.970 70.140 4.280 ;
        RECT 70.730 3.970 71.050 4.280 ;
        RECT 72.360 4.050 72.650 4.310 ;
        RECT 72.430 3.830 72.570 4.050 ;
        RECT 73.930 3.970 74.250 4.280 ;
        RECT 75.570 3.970 75.890 4.280 ;
        RECT 76.480 3.970 76.800 4.280 ;
        RECT 78.110 4.050 78.400 4.310 ;
        RECT 78.180 3.830 78.320 4.050 ;
        RECT 79.680 3.970 80.000 4.280 ;
        RECT 81.320 3.970 81.640 4.280 ;
        RECT 82.230 3.970 82.550 4.280 ;
        RECT 83.860 4.050 84.150 4.310 ;
        RECT 83.930 3.830 84.070 4.050 ;
        RECT 85.430 3.970 85.750 4.280 ;
        RECT 87.070 3.970 87.390 4.280 ;
        RECT 87.980 3.970 88.300 4.280 ;
        RECT 89.610 4.050 89.900 4.310 ;
        RECT 89.680 3.830 89.820 4.050 ;
        RECT 91.180 3.970 91.500 4.280 ;
        RECT 92.820 3.970 93.140 4.280 ;
        RECT 93.730 3.970 94.050 4.280 ;
        RECT 1.270 3.690 94.660 3.830 ;
        RECT 1.270 3.630 1.590 3.690 ;
        RECT 2.960 3.230 3.280 3.540 ;
        RECT 3.870 3.230 4.190 3.540 ;
        RECT 7.060 3.450 7.350 3.690 ;
        RECT 5.460 3.140 5.830 3.450 ;
        RECT 8.710 3.230 9.030 3.540 ;
        RECT 9.620 3.230 9.940 3.540 ;
        RECT 12.810 3.450 13.100 3.690 ;
        RECT 11.210 3.140 11.580 3.450 ;
        RECT 14.460 3.230 14.780 3.540 ;
        RECT 15.370 3.230 15.690 3.540 ;
        RECT 18.560 3.450 18.850 3.690 ;
        RECT 16.960 3.140 17.330 3.450 ;
        RECT 20.210 3.230 20.530 3.540 ;
        RECT 21.120 3.230 21.440 3.540 ;
        RECT 24.310 3.450 24.600 3.690 ;
        RECT 22.710 3.140 23.080 3.450 ;
        RECT 25.960 3.230 26.280 3.540 ;
        RECT 26.870 3.230 27.190 3.540 ;
        RECT 30.060 3.450 30.350 3.690 ;
        RECT 28.460 3.140 28.830 3.450 ;
        RECT 31.710 3.230 32.030 3.540 ;
        RECT 32.620 3.230 32.940 3.540 ;
        RECT 35.810 3.450 36.100 3.690 ;
        RECT 34.210 3.140 34.580 3.450 ;
        RECT 37.460 3.230 37.780 3.540 ;
        RECT 38.370 3.230 38.690 3.540 ;
        RECT 41.560 3.450 41.850 3.690 ;
        RECT 39.960 3.140 40.330 3.450 ;
        RECT 43.210 3.230 43.530 3.540 ;
        RECT 44.120 3.230 44.440 3.540 ;
        RECT 47.310 3.450 47.600 3.690 ;
        RECT 45.710 3.140 46.080 3.450 ;
        RECT 48.960 3.230 49.280 3.540 ;
        RECT 49.870 3.230 50.190 3.540 ;
        RECT 53.060 3.450 53.350 3.690 ;
        RECT 51.460 3.140 51.830 3.450 ;
        RECT 54.710 3.230 55.030 3.540 ;
        RECT 55.620 3.230 55.940 3.540 ;
        RECT 58.810 3.450 59.100 3.690 ;
        RECT 57.210 3.140 57.580 3.450 ;
        RECT 60.460 3.230 60.780 3.540 ;
        RECT 61.370 3.230 61.690 3.540 ;
        RECT 64.560 3.450 64.850 3.690 ;
        RECT 62.960 3.140 63.330 3.450 ;
        RECT 66.210 3.230 66.530 3.540 ;
        RECT 67.120 3.230 67.440 3.540 ;
        RECT 70.310 3.450 70.600 3.690 ;
        RECT 68.710 3.140 69.080 3.450 ;
        RECT 71.960 3.230 72.280 3.540 ;
        RECT 72.870 3.230 73.190 3.540 ;
        RECT 76.060 3.450 76.350 3.690 ;
        RECT 74.460 3.140 74.830 3.450 ;
        RECT 77.710 3.230 78.030 3.540 ;
        RECT 78.620 3.230 78.940 3.540 ;
        RECT 81.810 3.450 82.100 3.690 ;
        RECT 80.210 3.140 80.580 3.450 ;
        RECT 83.460 3.230 83.780 3.540 ;
        RECT 84.370 3.230 84.690 3.540 ;
        RECT 87.560 3.450 87.850 3.690 ;
        RECT 85.960 3.140 86.330 3.450 ;
        RECT 89.210 3.230 89.530 3.540 ;
        RECT 90.120 3.230 90.440 3.540 ;
        RECT 93.310 3.450 93.600 3.690 ;
        RECT 91.710 3.140 92.080 3.450 ;
        RECT 3.360 1.640 3.650 1.900 ;
        RECT 1.260 1.420 1.580 1.480 ;
        RECT 3.430 1.420 3.570 1.640 ;
        RECT 4.930 1.560 5.250 1.870 ;
        RECT 6.570 1.560 6.890 1.870 ;
        RECT 7.480 1.560 7.800 1.870 ;
        RECT 9.110 1.640 9.400 1.900 ;
        RECT 9.180 1.420 9.320 1.640 ;
        RECT 10.680 1.560 11.000 1.870 ;
        RECT 12.320 1.560 12.640 1.870 ;
        RECT 13.230 1.560 13.550 1.870 ;
        RECT 14.860 1.640 15.150 1.900 ;
        RECT 14.930 1.420 15.070 1.640 ;
        RECT 16.430 1.560 16.750 1.870 ;
        RECT 18.070 1.560 18.390 1.870 ;
        RECT 18.980 1.560 19.300 1.870 ;
        RECT 20.610 1.640 20.900 1.900 ;
        RECT 20.680 1.420 20.820 1.640 ;
        RECT 22.180 1.560 22.500 1.870 ;
        RECT 23.820 1.560 24.140 1.870 ;
        RECT 24.730 1.560 25.050 1.870 ;
        RECT 26.360 1.640 26.650 1.900 ;
        RECT 26.430 1.420 26.570 1.640 ;
        RECT 27.930 1.560 28.250 1.870 ;
        RECT 29.570 1.560 29.890 1.870 ;
        RECT 30.480 1.560 30.800 1.870 ;
        RECT 32.110 1.640 32.400 1.900 ;
        RECT 32.180 1.420 32.320 1.640 ;
        RECT 33.680 1.560 34.000 1.870 ;
        RECT 35.320 1.560 35.640 1.870 ;
        RECT 36.230 1.560 36.550 1.870 ;
        RECT 37.860 1.640 38.150 1.900 ;
        RECT 37.930 1.420 38.070 1.640 ;
        RECT 39.430 1.560 39.750 1.870 ;
        RECT 41.070 1.560 41.390 1.870 ;
        RECT 41.980 1.560 42.300 1.870 ;
        RECT 43.610 1.640 43.900 1.900 ;
        RECT 43.680 1.420 43.820 1.640 ;
        RECT 45.180 1.560 45.500 1.870 ;
        RECT 46.820 1.560 47.140 1.870 ;
        RECT 47.730 1.560 48.050 1.870 ;
        RECT 49.360 1.640 49.650 1.900 ;
        RECT 49.430 1.420 49.570 1.640 ;
        RECT 50.930 1.560 51.250 1.870 ;
        RECT 52.570 1.560 52.890 1.870 ;
        RECT 53.480 1.560 53.800 1.870 ;
        RECT 55.110 1.640 55.400 1.900 ;
        RECT 55.180 1.420 55.320 1.640 ;
        RECT 56.680 1.560 57.000 1.870 ;
        RECT 58.320 1.560 58.640 1.870 ;
        RECT 59.230 1.560 59.550 1.870 ;
        RECT 60.860 1.640 61.150 1.900 ;
        RECT 60.930 1.420 61.070 1.640 ;
        RECT 62.430 1.560 62.750 1.870 ;
        RECT 64.070 1.560 64.390 1.870 ;
        RECT 64.980 1.560 65.300 1.870 ;
        RECT 66.610 1.640 66.900 1.900 ;
        RECT 66.680 1.420 66.820 1.640 ;
        RECT 68.180 1.560 68.500 1.870 ;
        RECT 69.820 1.560 70.140 1.870 ;
        RECT 70.730 1.560 71.050 1.870 ;
        RECT 72.360 1.640 72.650 1.900 ;
        RECT 72.430 1.420 72.570 1.640 ;
        RECT 73.930 1.560 74.250 1.870 ;
        RECT 75.570 1.560 75.890 1.870 ;
        RECT 76.480 1.560 76.800 1.870 ;
        RECT 78.110 1.640 78.400 1.900 ;
        RECT 78.180 1.420 78.320 1.640 ;
        RECT 79.680 1.560 80.000 1.870 ;
        RECT 81.320 1.560 81.640 1.870 ;
        RECT 82.230 1.560 82.550 1.870 ;
        RECT 83.860 1.640 84.150 1.900 ;
        RECT 83.930 1.420 84.070 1.640 ;
        RECT 85.430 1.560 85.750 1.870 ;
        RECT 87.070 1.560 87.390 1.870 ;
        RECT 87.980 1.560 88.300 1.870 ;
        RECT 89.610 1.640 89.900 1.900 ;
        RECT 89.680 1.420 89.820 1.640 ;
        RECT 91.180 1.560 91.500 1.870 ;
        RECT 92.820 1.560 93.140 1.870 ;
        RECT 93.730 1.560 94.050 1.870 ;
        RECT 1.260 1.280 94.660 1.420 ;
        RECT 1.260 1.220 1.580 1.280 ;
        RECT 2.960 0.820 3.280 1.130 ;
        RECT 3.870 0.820 4.190 1.130 ;
        RECT 7.060 1.040 7.350 1.280 ;
        RECT 5.460 0.730 5.830 1.040 ;
        RECT 8.710 0.820 9.030 1.130 ;
        RECT 9.620 0.820 9.940 1.130 ;
        RECT 12.810 1.040 13.100 1.280 ;
        RECT 11.210 0.730 11.580 1.040 ;
        RECT 14.460 0.820 14.780 1.130 ;
        RECT 15.370 0.820 15.690 1.130 ;
        RECT 18.560 1.040 18.850 1.280 ;
        RECT 16.960 0.730 17.330 1.040 ;
        RECT 20.210 0.820 20.530 1.130 ;
        RECT 21.120 0.820 21.440 1.130 ;
        RECT 24.310 1.040 24.600 1.280 ;
        RECT 22.710 0.730 23.080 1.040 ;
        RECT 25.960 0.820 26.280 1.130 ;
        RECT 26.870 0.820 27.190 1.130 ;
        RECT 30.060 1.040 30.350 1.280 ;
        RECT 28.460 0.730 28.830 1.040 ;
        RECT 31.710 0.820 32.030 1.130 ;
        RECT 32.620 0.820 32.940 1.130 ;
        RECT 35.810 1.040 36.100 1.280 ;
        RECT 34.210 0.730 34.580 1.040 ;
        RECT 37.460 0.820 37.780 1.130 ;
        RECT 38.370 0.820 38.690 1.130 ;
        RECT 41.560 1.040 41.850 1.280 ;
        RECT 39.960 0.730 40.330 1.040 ;
        RECT 43.210 0.820 43.530 1.130 ;
        RECT 44.120 0.820 44.440 1.130 ;
        RECT 47.310 1.040 47.600 1.280 ;
        RECT 45.710 0.730 46.080 1.040 ;
        RECT 48.960 0.820 49.280 1.130 ;
        RECT 49.870 0.820 50.190 1.130 ;
        RECT 53.060 1.040 53.350 1.280 ;
        RECT 51.460 0.730 51.830 1.040 ;
        RECT 54.710 0.820 55.030 1.130 ;
        RECT 55.620 0.820 55.940 1.130 ;
        RECT 58.810 1.040 59.100 1.280 ;
        RECT 57.210 0.730 57.580 1.040 ;
        RECT 60.460 0.820 60.780 1.130 ;
        RECT 61.370 0.820 61.690 1.130 ;
        RECT 64.560 1.040 64.850 1.280 ;
        RECT 62.960 0.730 63.330 1.040 ;
        RECT 66.210 0.820 66.530 1.130 ;
        RECT 67.120 0.820 67.440 1.130 ;
        RECT 70.310 1.040 70.600 1.280 ;
        RECT 68.710 0.730 69.080 1.040 ;
        RECT 71.960 0.820 72.280 1.130 ;
        RECT 72.870 0.820 73.190 1.130 ;
        RECT 76.060 1.040 76.350 1.280 ;
        RECT 74.460 0.730 74.830 1.040 ;
        RECT 77.710 0.820 78.030 1.130 ;
        RECT 78.620 0.820 78.940 1.130 ;
        RECT 81.810 1.040 82.100 1.280 ;
        RECT 80.210 0.730 80.580 1.040 ;
        RECT 83.460 0.820 83.780 1.130 ;
        RECT 84.370 0.820 84.690 1.130 ;
        RECT 87.560 1.040 87.850 1.280 ;
        RECT 85.960 0.730 86.330 1.040 ;
        RECT 89.210 0.820 89.530 1.130 ;
        RECT 90.120 0.820 90.440 1.130 ;
        RECT 93.310 1.040 93.600 1.280 ;
        RECT 91.710 0.730 92.080 1.040 ;
        RECT 3.360 -0.770 3.650 -0.510 ;
        RECT 1.260 -0.990 1.580 -0.900 ;
        RECT 3.430 -0.990 3.570 -0.770 ;
        RECT 4.930 -0.850 5.250 -0.540 ;
        RECT 6.570 -0.850 6.890 -0.540 ;
        RECT 7.480 -0.850 7.800 -0.540 ;
        RECT 9.110 -0.770 9.400 -0.510 ;
        RECT 9.180 -0.990 9.320 -0.770 ;
        RECT 10.680 -0.850 11.000 -0.540 ;
        RECT 12.320 -0.850 12.640 -0.540 ;
        RECT 13.230 -0.850 13.550 -0.540 ;
        RECT 14.860 -0.770 15.150 -0.510 ;
        RECT 14.930 -0.990 15.070 -0.770 ;
        RECT 16.430 -0.850 16.750 -0.540 ;
        RECT 18.070 -0.850 18.390 -0.540 ;
        RECT 18.980 -0.850 19.300 -0.540 ;
        RECT 20.610 -0.770 20.900 -0.510 ;
        RECT 20.680 -0.990 20.820 -0.770 ;
        RECT 22.180 -0.850 22.500 -0.540 ;
        RECT 23.820 -0.850 24.140 -0.540 ;
        RECT 24.730 -0.850 25.050 -0.540 ;
        RECT 26.360 -0.770 26.650 -0.510 ;
        RECT 26.430 -0.990 26.570 -0.770 ;
        RECT 27.930 -0.850 28.250 -0.540 ;
        RECT 29.570 -0.850 29.890 -0.540 ;
        RECT 30.480 -0.850 30.800 -0.540 ;
        RECT 32.110 -0.770 32.400 -0.510 ;
        RECT 32.180 -0.990 32.320 -0.770 ;
        RECT 33.680 -0.850 34.000 -0.540 ;
        RECT 35.320 -0.850 35.640 -0.540 ;
        RECT 36.230 -0.850 36.550 -0.540 ;
        RECT 37.860 -0.770 38.150 -0.510 ;
        RECT 37.930 -0.990 38.070 -0.770 ;
        RECT 39.430 -0.850 39.750 -0.540 ;
        RECT 41.070 -0.850 41.390 -0.540 ;
        RECT 41.980 -0.850 42.300 -0.540 ;
        RECT 43.610 -0.770 43.900 -0.510 ;
        RECT 43.680 -0.990 43.820 -0.770 ;
        RECT 45.180 -0.850 45.500 -0.540 ;
        RECT 46.820 -0.850 47.140 -0.540 ;
        RECT 47.730 -0.850 48.050 -0.540 ;
        RECT 49.360 -0.770 49.650 -0.510 ;
        RECT 49.430 -0.990 49.570 -0.770 ;
        RECT 50.930 -0.850 51.250 -0.540 ;
        RECT 52.570 -0.850 52.890 -0.540 ;
        RECT 53.480 -0.850 53.800 -0.540 ;
        RECT 55.110 -0.770 55.400 -0.510 ;
        RECT 55.180 -0.990 55.320 -0.770 ;
        RECT 56.680 -0.850 57.000 -0.540 ;
        RECT 58.320 -0.850 58.640 -0.540 ;
        RECT 59.230 -0.850 59.550 -0.540 ;
        RECT 60.860 -0.770 61.150 -0.510 ;
        RECT 60.930 -0.990 61.070 -0.770 ;
        RECT 62.430 -0.850 62.750 -0.540 ;
        RECT 64.070 -0.850 64.390 -0.540 ;
        RECT 64.980 -0.850 65.300 -0.540 ;
        RECT 66.610 -0.770 66.900 -0.510 ;
        RECT 66.680 -0.990 66.820 -0.770 ;
        RECT 68.180 -0.850 68.500 -0.540 ;
        RECT 69.820 -0.850 70.140 -0.540 ;
        RECT 70.730 -0.850 71.050 -0.540 ;
        RECT 72.360 -0.770 72.650 -0.510 ;
        RECT 72.430 -0.990 72.570 -0.770 ;
        RECT 73.930 -0.850 74.250 -0.540 ;
        RECT 75.570 -0.850 75.890 -0.540 ;
        RECT 76.480 -0.850 76.800 -0.540 ;
        RECT 78.110 -0.770 78.400 -0.510 ;
        RECT 78.180 -0.990 78.320 -0.770 ;
        RECT 79.680 -0.850 80.000 -0.540 ;
        RECT 81.320 -0.850 81.640 -0.540 ;
        RECT 82.230 -0.850 82.550 -0.540 ;
        RECT 83.860 -0.770 84.150 -0.510 ;
        RECT 83.930 -0.990 84.070 -0.770 ;
        RECT 85.430 -0.850 85.750 -0.540 ;
        RECT 87.070 -0.850 87.390 -0.540 ;
        RECT 87.980 -0.850 88.300 -0.540 ;
        RECT 89.610 -0.770 89.900 -0.510 ;
        RECT 89.680 -0.990 89.820 -0.770 ;
        RECT 91.180 -0.850 91.500 -0.540 ;
        RECT 92.820 -0.850 93.140 -0.540 ;
        RECT 93.730 -0.850 94.050 -0.540 ;
        RECT 1.260 -1.130 94.660 -0.990 ;
        RECT 1.260 -1.220 1.580 -1.130 ;
        RECT 2.960 -1.590 3.280 -1.280 ;
        RECT 3.870 -1.590 4.190 -1.280 ;
        RECT 7.060 -1.370 7.350 -1.130 ;
        RECT 5.460 -1.680 5.830 -1.370 ;
        RECT 8.710 -1.590 9.030 -1.280 ;
        RECT 9.620 -1.590 9.940 -1.280 ;
        RECT 12.810 -1.370 13.100 -1.130 ;
        RECT 11.210 -1.680 11.580 -1.370 ;
        RECT 14.460 -1.590 14.780 -1.280 ;
        RECT 15.370 -1.590 15.690 -1.280 ;
        RECT 18.560 -1.370 18.850 -1.130 ;
        RECT 16.960 -1.680 17.330 -1.370 ;
        RECT 20.210 -1.590 20.530 -1.280 ;
        RECT 21.120 -1.590 21.440 -1.280 ;
        RECT 24.310 -1.370 24.600 -1.130 ;
        RECT 22.710 -1.680 23.080 -1.370 ;
        RECT 25.960 -1.590 26.280 -1.280 ;
        RECT 26.870 -1.590 27.190 -1.280 ;
        RECT 30.060 -1.370 30.350 -1.130 ;
        RECT 28.460 -1.680 28.830 -1.370 ;
        RECT 31.710 -1.590 32.030 -1.280 ;
        RECT 32.620 -1.590 32.940 -1.280 ;
        RECT 35.810 -1.370 36.100 -1.130 ;
        RECT 34.210 -1.680 34.580 -1.370 ;
        RECT 37.460 -1.590 37.780 -1.280 ;
        RECT 38.370 -1.590 38.690 -1.280 ;
        RECT 41.560 -1.370 41.850 -1.130 ;
        RECT 39.960 -1.680 40.330 -1.370 ;
        RECT 43.210 -1.590 43.530 -1.280 ;
        RECT 44.120 -1.590 44.440 -1.280 ;
        RECT 47.310 -1.370 47.600 -1.130 ;
        RECT 45.710 -1.680 46.080 -1.370 ;
        RECT 48.960 -1.590 49.280 -1.280 ;
        RECT 49.870 -1.590 50.190 -1.280 ;
        RECT 53.060 -1.370 53.350 -1.130 ;
        RECT 51.460 -1.680 51.830 -1.370 ;
        RECT 54.710 -1.590 55.030 -1.280 ;
        RECT 55.620 -1.590 55.940 -1.280 ;
        RECT 58.810 -1.370 59.100 -1.130 ;
        RECT 57.210 -1.680 57.580 -1.370 ;
        RECT 60.460 -1.590 60.780 -1.280 ;
        RECT 61.370 -1.590 61.690 -1.280 ;
        RECT 64.560 -1.370 64.850 -1.130 ;
        RECT 62.960 -1.680 63.330 -1.370 ;
        RECT 66.210 -1.590 66.530 -1.280 ;
        RECT 67.120 -1.590 67.440 -1.280 ;
        RECT 70.310 -1.370 70.600 -1.130 ;
        RECT 68.710 -1.680 69.080 -1.370 ;
        RECT 71.960 -1.590 72.280 -1.280 ;
        RECT 72.870 -1.590 73.190 -1.280 ;
        RECT 76.060 -1.370 76.350 -1.130 ;
        RECT 74.460 -1.680 74.830 -1.370 ;
        RECT 77.710 -1.590 78.030 -1.280 ;
        RECT 78.620 -1.590 78.940 -1.280 ;
        RECT 81.810 -1.370 82.100 -1.130 ;
        RECT 80.210 -1.680 80.580 -1.370 ;
        RECT 83.460 -1.590 83.780 -1.280 ;
        RECT 84.370 -1.590 84.690 -1.280 ;
        RECT 87.560 -1.370 87.850 -1.130 ;
        RECT 85.960 -1.680 86.330 -1.370 ;
        RECT 89.210 -1.590 89.530 -1.280 ;
        RECT 90.120 -1.590 90.440 -1.280 ;
        RECT 93.310 -1.370 93.600 -1.130 ;
        RECT 91.710 -1.680 92.080 -1.370 ;
        RECT 1.260 -1.820 1.580 -1.750 ;
        RECT 2.460 -1.820 2.760 -1.750 ;
        RECT 8.210 -1.820 8.510 -1.750 ;
        RECT 13.960 -1.820 14.260 -1.750 ;
        RECT 19.710 -1.820 20.010 -1.750 ;
        RECT 25.460 -1.820 25.760 -1.750 ;
        RECT 31.210 -1.820 31.510 -1.750 ;
        RECT 36.960 -1.820 37.260 -1.750 ;
        RECT 42.710 -1.820 43.010 -1.750 ;
        RECT 48.460 -1.820 48.760 -1.750 ;
        RECT 54.210 -1.820 54.510 -1.750 ;
        RECT 59.960 -1.820 60.260 -1.750 ;
        RECT 65.710 -1.820 66.010 -1.750 ;
        RECT 71.460 -1.820 71.760 -1.750 ;
        RECT 77.210 -1.820 77.510 -1.750 ;
        RECT 82.960 -1.820 83.260 -1.750 ;
        RECT 88.710 -1.820 89.010 -1.750 ;
        RECT 1.260 -1.960 94.660 -1.820 ;
        RECT 1.260 -2.070 1.580 -1.960 ;
        RECT 2.460 -2.040 2.760 -1.960 ;
        RECT 8.210 -2.040 8.510 -1.960 ;
        RECT 13.960 -2.040 14.260 -1.960 ;
        RECT 19.710 -2.040 20.010 -1.960 ;
        RECT 25.460 -2.040 25.760 -1.960 ;
        RECT 31.210 -2.040 31.510 -1.960 ;
        RECT 36.960 -2.040 37.260 -1.960 ;
        RECT 42.710 -2.040 43.010 -1.960 ;
        RECT 48.460 -2.040 48.760 -1.960 ;
        RECT 54.210 -2.040 54.510 -1.960 ;
        RECT 59.960 -2.040 60.260 -1.960 ;
        RECT 65.710 -2.040 66.010 -1.960 ;
        RECT 71.460 -2.040 71.760 -1.960 ;
        RECT 77.210 -2.040 77.510 -1.960 ;
        RECT 82.960 -2.040 83.260 -1.960 ;
        RECT 88.710 -2.040 89.010 -1.960 ;
        RECT 1.260 -2.630 1.580 -2.540 ;
        RECT 8.010 -2.630 8.310 -2.530 ;
        RECT 13.760 -2.630 14.060 -2.530 ;
        RECT 19.510 -2.630 19.810 -2.530 ;
        RECT 25.260 -2.630 25.560 -2.530 ;
        RECT 31.010 -2.630 31.310 -2.530 ;
        RECT 36.760 -2.630 37.060 -2.530 ;
        RECT 42.510 -2.630 42.810 -2.530 ;
        RECT 48.260 -2.630 48.560 -2.530 ;
        RECT 54.010 -2.630 54.310 -2.530 ;
        RECT 59.760 -2.630 60.060 -2.530 ;
        RECT 65.510 -2.630 65.810 -2.530 ;
        RECT 71.260 -2.630 71.560 -2.530 ;
        RECT 77.010 -2.630 77.310 -2.530 ;
        RECT 82.760 -2.630 83.060 -2.530 ;
        RECT 88.510 -2.630 88.810 -2.530 ;
        RECT 94.260 -2.630 94.560 -2.530 ;
        RECT 1.260 -2.770 94.660 -2.630 ;
        RECT 1.260 -2.860 1.580 -2.770 ;
        RECT 8.010 -2.860 8.310 -2.770 ;
        RECT 13.760 -2.860 14.060 -2.770 ;
        RECT 19.510 -2.860 19.810 -2.770 ;
        RECT 25.260 -2.860 25.560 -2.770 ;
        RECT 31.010 -2.860 31.310 -2.770 ;
        RECT 36.760 -2.860 37.060 -2.770 ;
        RECT 42.510 -2.860 42.810 -2.770 ;
        RECT 48.260 -2.860 48.560 -2.770 ;
        RECT 54.010 -2.860 54.310 -2.770 ;
        RECT 59.760 -2.860 60.060 -2.770 ;
        RECT 65.510 -2.860 65.810 -2.770 ;
        RECT 71.260 -2.860 71.560 -2.770 ;
        RECT 77.010 -2.860 77.310 -2.770 ;
        RECT 82.760 -2.860 83.060 -2.770 ;
        RECT 88.510 -2.860 88.810 -2.770 ;
        RECT 94.260 -2.860 94.560 -2.770 ;
        RECT 3.360 -3.180 3.650 -2.920 ;
        RECT 1.290 -3.400 1.550 -3.310 ;
        RECT 3.430 -3.400 3.570 -3.180 ;
        RECT 4.930 -3.260 5.250 -2.950 ;
        RECT 6.570 -3.260 6.890 -2.950 ;
        RECT 7.480 -3.260 7.800 -2.950 ;
        RECT 9.110 -3.180 9.400 -2.920 ;
        RECT 9.180 -3.400 9.320 -3.180 ;
        RECT 10.680 -3.260 11.000 -2.950 ;
        RECT 12.320 -3.260 12.640 -2.950 ;
        RECT 13.230 -3.260 13.550 -2.950 ;
        RECT 14.860 -3.180 15.150 -2.920 ;
        RECT 14.930 -3.400 15.070 -3.180 ;
        RECT 16.430 -3.260 16.750 -2.950 ;
        RECT 18.070 -3.260 18.390 -2.950 ;
        RECT 18.980 -3.260 19.300 -2.950 ;
        RECT 20.610 -3.180 20.900 -2.920 ;
        RECT 20.680 -3.400 20.820 -3.180 ;
        RECT 22.180 -3.260 22.500 -2.950 ;
        RECT 23.820 -3.260 24.140 -2.950 ;
        RECT 24.730 -3.260 25.050 -2.950 ;
        RECT 26.360 -3.180 26.650 -2.920 ;
        RECT 26.430 -3.400 26.570 -3.180 ;
        RECT 27.930 -3.260 28.250 -2.950 ;
        RECT 29.570 -3.260 29.890 -2.950 ;
        RECT 30.480 -3.260 30.800 -2.950 ;
        RECT 32.110 -3.180 32.400 -2.920 ;
        RECT 32.180 -3.400 32.320 -3.180 ;
        RECT 33.680 -3.260 34.000 -2.950 ;
        RECT 35.320 -3.260 35.640 -2.950 ;
        RECT 36.230 -3.260 36.550 -2.950 ;
        RECT 37.860 -3.180 38.150 -2.920 ;
        RECT 37.930 -3.400 38.070 -3.180 ;
        RECT 39.430 -3.260 39.750 -2.950 ;
        RECT 41.070 -3.260 41.390 -2.950 ;
        RECT 41.980 -3.260 42.300 -2.950 ;
        RECT 43.610 -3.180 43.900 -2.920 ;
        RECT 43.680 -3.400 43.820 -3.180 ;
        RECT 45.180 -3.260 45.500 -2.950 ;
        RECT 46.820 -3.260 47.140 -2.950 ;
        RECT 47.730 -3.260 48.050 -2.950 ;
        RECT 49.360 -3.180 49.650 -2.920 ;
        RECT 49.430 -3.400 49.570 -3.180 ;
        RECT 50.930 -3.260 51.250 -2.950 ;
        RECT 52.570 -3.260 52.890 -2.950 ;
        RECT 53.480 -3.260 53.800 -2.950 ;
        RECT 55.110 -3.180 55.400 -2.920 ;
        RECT 55.180 -3.400 55.320 -3.180 ;
        RECT 56.680 -3.260 57.000 -2.950 ;
        RECT 58.320 -3.260 58.640 -2.950 ;
        RECT 59.230 -3.260 59.550 -2.950 ;
        RECT 60.860 -3.180 61.150 -2.920 ;
        RECT 60.930 -3.400 61.070 -3.180 ;
        RECT 62.430 -3.260 62.750 -2.950 ;
        RECT 64.070 -3.260 64.390 -2.950 ;
        RECT 64.980 -3.260 65.300 -2.950 ;
        RECT 66.610 -3.180 66.900 -2.920 ;
        RECT 66.680 -3.400 66.820 -3.180 ;
        RECT 68.180 -3.260 68.500 -2.950 ;
        RECT 69.820 -3.260 70.140 -2.950 ;
        RECT 70.730 -3.260 71.050 -2.950 ;
        RECT 72.360 -3.180 72.650 -2.920 ;
        RECT 72.430 -3.400 72.570 -3.180 ;
        RECT 73.930 -3.260 74.250 -2.950 ;
        RECT 75.570 -3.260 75.890 -2.950 ;
        RECT 76.480 -3.260 76.800 -2.950 ;
        RECT 78.110 -3.180 78.400 -2.920 ;
        RECT 78.180 -3.400 78.320 -3.180 ;
        RECT 79.680 -3.260 80.000 -2.950 ;
        RECT 81.320 -3.260 81.640 -2.950 ;
        RECT 82.230 -3.260 82.550 -2.950 ;
        RECT 83.860 -3.180 84.150 -2.920 ;
        RECT 83.930 -3.400 84.070 -3.180 ;
        RECT 85.430 -3.260 85.750 -2.950 ;
        RECT 87.070 -3.260 87.390 -2.950 ;
        RECT 87.980 -3.260 88.300 -2.950 ;
        RECT 89.610 -3.180 89.900 -2.920 ;
        RECT 89.680 -3.400 89.820 -3.180 ;
        RECT 91.180 -3.260 91.500 -2.950 ;
        RECT 92.820 -3.260 93.140 -2.950 ;
        RECT 93.730 -3.260 94.050 -2.950 ;
        RECT 1.290 -3.540 94.660 -3.400 ;
        RECT 1.290 -3.630 1.550 -3.540 ;
        RECT 2.960 -4.000 3.280 -3.690 ;
        RECT 3.870 -4.000 4.190 -3.690 ;
        RECT 7.060 -3.780 7.350 -3.540 ;
        RECT 5.460 -4.090 5.830 -3.780 ;
        RECT 8.710 -4.000 9.030 -3.690 ;
        RECT 9.620 -4.000 9.940 -3.690 ;
        RECT 12.810 -3.780 13.100 -3.540 ;
        RECT 11.210 -4.090 11.580 -3.780 ;
        RECT 14.460 -4.000 14.780 -3.690 ;
        RECT 15.370 -4.000 15.690 -3.690 ;
        RECT 18.560 -3.780 18.850 -3.540 ;
        RECT 16.960 -4.090 17.330 -3.780 ;
        RECT 20.210 -4.000 20.530 -3.690 ;
        RECT 21.120 -4.000 21.440 -3.690 ;
        RECT 24.310 -3.780 24.600 -3.540 ;
        RECT 22.710 -4.090 23.080 -3.780 ;
        RECT 25.960 -4.000 26.280 -3.690 ;
        RECT 26.870 -4.000 27.190 -3.690 ;
        RECT 30.060 -3.780 30.350 -3.540 ;
        RECT 28.460 -4.090 28.830 -3.780 ;
        RECT 31.710 -4.000 32.030 -3.690 ;
        RECT 32.620 -4.000 32.940 -3.690 ;
        RECT 35.810 -3.780 36.100 -3.540 ;
        RECT 34.210 -4.090 34.580 -3.780 ;
        RECT 37.460 -4.000 37.780 -3.690 ;
        RECT 38.370 -4.000 38.690 -3.690 ;
        RECT 41.560 -3.780 41.850 -3.540 ;
        RECT 39.960 -4.090 40.330 -3.780 ;
        RECT 43.210 -4.000 43.530 -3.690 ;
        RECT 44.120 -4.000 44.440 -3.690 ;
        RECT 47.310 -3.780 47.600 -3.540 ;
        RECT 45.710 -4.090 46.080 -3.780 ;
        RECT 48.960 -4.000 49.280 -3.690 ;
        RECT 49.870 -4.000 50.190 -3.690 ;
        RECT 53.060 -3.780 53.350 -3.540 ;
        RECT 51.460 -4.090 51.830 -3.780 ;
        RECT 54.710 -4.000 55.030 -3.690 ;
        RECT 55.620 -4.000 55.940 -3.690 ;
        RECT 58.810 -3.780 59.100 -3.540 ;
        RECT 57.210 -4.090 57.580 -3.780 ;
        RECT 60.460 -4.000 60.780 -3.690 ;
        RECT 61.370 -4.000 61.690 -3.690 ;
        RECT 64.560 -3.780 64.850 -3.540 ;
        RECT 62.960 -4.090 63.330 -3.780 ;
        RECT 66.210 -4.000 66.530 -3.690 ;
        RECT 67.120 -4.000 67.440 -3.690 ;
        RECT 70.310 -3.780 70.600 -3.540 ;
        RECT 68.710 -4.090 69.080 -3.780 ;
        RECT 71.960 -4.000 72.280 -3.690 ;
        RECT 72.870 -4.000 73.190 -3.690 ;
        RECT 76.060 -3.780 76.350 -3.540 ;
        RECT 74.460 -4.090 74.830 -3.780 ;
        RECT 77.710 -4.000 78.030 -3.690 ;
        RECT 78.620 -4.000 78.940 -3.690 ;
        RECT 81.810 -3.780 82.100 -3.540 ;
        RECT 80.210 -4.090 80.580 -3.780 ;
        RECT 83.460 -4.000 83.780 -3.690 ;
        RECT 84.370 -4.000 84.690 -3.690 ;
        RECT 87.560 -3.780 87.850 -3.540 ;
        RECT 85.960 -4.090 86.330 -3.780 ;
        RECT 89.210 -4.000 89.530 -3.690 ;
        RECT 90.120 -4.000 90.440 -3.690 ;
        RECT 93.310 -3.780 93.600 -3.540 ;
        RECT 91.710 -4.090 92.080 -3.780 ;
        RECT 1.260 -4.230 1.580 -4.130 ;
        RECT 2.460 -4.230 2.760 -4.160 ;
        RECT 8.210 -4.230 8.510 -4.160 ;
        RECT 13.960 -4.230 14.260 -4.160 ;
        RECT 19.710 -4.230 20.010 -4.160 ;
        RECT 25.460 -4.230 25.760 -4.160 ;
        RECT 31.210 -4.230 31.510 -4.160 ;
        RECT 36.960 -4.230 37.260 -4.160 ;
        RECT 42.710 -4.230 43.010 -4.160 ;
        RECT 48.460 -4.230 48.760 -4.160 ;
        RECT 54.210 -4.230 54.510 -4.160 ;
        RECT 59.960 -4.230 60.260 -4.160 ;
        RECT 65.710 -4.230 66.010 -4.160 ;
        RECT 71.460 -4.230 71.760 -4.160 ;
        RECT 77.210 -4.230 77.510 -4.160 ;
        RECT 82.960 -4.230 83.260 -4.160 ;
        RECT 88.710 -4.230 89.010 -4.160 ;
        RECT 1.260 -4.370 94.660 -4.230 ;
        RECT 1.260 -4.450 1.580 -4.370 ;
        RECT 2.460 -4.450 2.760 -4.370 ;
        RECT 8.210 -4.450 8.510 -4.370 ;
        RECT 13.960 -4.450 14.260 -4.370 ;
        RECT 19.710 -4.450 20.010 -4.370 ;
        RECT 25.460 -4.450 25.760 -4.370 ;
        RECT 31.210 -4.450 31.510 -4.370 ;
        RECT 36.960 -4.450 37.260 -4.370 ;
        RECT 42.710 -4.450 43.010 -4.370 ;
        RECT 48.460 -4.450 48.760 -4.370 ;
        RECT 54.210 -4.450 54.510 -4.370 ;
        RECT 59.960 -4.450 60.260 -4.370 ;
        RECT 65.710 -4.450 66.010 -4.370 ;
        RECT 71.460 -4.450 71.760 -4.370 ;
        RECT 77.210 -4.450 77.510 -4.370 ;
        RECT 82.960 -4.450 83.260 -4.370 ;
        RECT 88.710 -4.450 89.010 -4.370 ;
        RECT 1.270 -5.040 1.590 -4.920 ;
        RECT 8.010 -5.040 8.310 -4.940 ;
        RECT 13.760 -5.040 14.060 -4.940 ;
        RECT 19.510 -5.040 19.810 -4.940 ;
        RECT 25.260 -5.040 25.560 -4.940 ;
        RECT 31.010 -5.040 31.310 -4.940 ;
        RECT 36.760 -5.040 37.060 -4.940 ;
        RECT 42.510 -5.040 42.810 -4.940 ;
        RECT 48.260 -5.040 48.560 -4.940 ;
        RECT 54.010 -5.040 54.310 -4.940 ;
        RECT 59.760 -5.040 60.060 -4.940 ;
        RECT 65.510 -5.040 65.810 -4.940 ;
        RECT 71.260 -5.040 71.560 -4.940 ;
        RECT 77.010 -5.040 77.310 -4.940 ;
        RECT 82.760 -5.040 83.060 -4.940 ;
        RECT 88.510 -5.040 88.810 -4.940 ;
        RECT 94.260 -5.040 94.560 -4.940 ;
        RECT 1.270 -5.180 94.660 -5.040 ;
        RECT 1.270 -5.240 1.590 -5.180 ;
        RECT 8.010 -5.270 8.310 -5.180 ;
        RECT 13.760 -5.270 14.060 -5.180 ;
        RECT 19.510 -5.270 19.810 -5.180 ;
        RECT 25.260 -5.270 25.560 -5.180 ;
        RECT 31.010 -5.270 31.310 -5.180 ;
        RECT 36.760 -5.270 37.060 -5.180 ;
        RECT 42.510 -5.270 42.810 -5.180 ;
        RECT 48.260 -5.270 48.560 -5.180 ;
        RECT 54.010 -5.270 54.310 -5.180 ;
        RECT 59.760 -5.270 60.060 -5.180 ;
        RECT 65.510 -5.270 65.810 -5.180 ;
        RECT 71.260 -5.270 71.560 -5.180 ;
        RECT 77.010 -5.270 77.310 -5.180 ;
        RECT 82.760 -5.270 83.060 -5.180 ;
        RECT 88.510 -5.270 88.810 -5.180 ;
        RECT 94.260 -5.270 94.560 -5.180 ;
        RECT 3.360 -5.590 3.650 -5.330 ;
        RECT 1.260 -5.810 1.580 -5.750 ;
        RECT 3.430 -5.810 3.570 -5.590 ;
        RECT 4.930 -5.670 5.250 -5.360 ;
        RECT 6.570 -5.670 6.890 -5.360 ;
        RECT 7.480 -5.670 7.800 -5.360 ;
        RECT 9.110 -5.590 9.400 -5.330 ;
        RECT 9.180 -5.810 9.320 -5.590 ;
        RECT 10.680 -5.670 11.000 -5.360 ;
        RECT 12.320 -5.670 12.640 -5.360 ;
        RECT 13.230 -5.670 13.550 -5.360 ;
        RECT 14.860 -5.590 15.150 -5.330 ;
        RECT 14.930 -5.810 15.070 -5.590 ;
        RECT 16.430 -5.670 16.750 -5.360 ;
        RECT 18.070 -5.670 18.390 -5.360 ;
        RECT 18.980 -5.670 19.300 -5.360 ;
        RECT 20.610 -5.590 20.900 -5.330 ;
        RECT 20.680 -5.810 20.820 -5.590 ;
        RECT 22.180 -5.670 22.500 -5.360 ;
        RECT 23.820 -5.670 24.140 -5.360 ;
        RECT 24.730 -5.670 25.050 -5.360 ;
        RECT 26.360 -5.590 26.650 -5.330 ;
        RECT 26.430 -5.810 26.570 -5.590 ;
        RECT 27.930 -5.670 28.250 -5.360 ;
        RECT 29.570 -5.670 29.890 -5.360 ;
        RECT 30.480 -5.670 30.800 -5.360 ;
        RECT 32.110 -5.590 32.400 -5.330 ;
        RECT 32.180 -5.810 32.320 -5.590 ;
        RECT 33.680 -5.670 34.000 -5.360 ;
        RECT 35.320 -5.670 35.640 -5.360 ;
        RECT 36.230 -5.670 36.550 -5.360 ;
        RECT 37.860 -5.590 38.150 -5.330 ;
        RECT 37.930 -5.810 38.070 -5.590 ;
        RECT 39.430 -5.670 39.750 -5.360 ;
        RECT 41.070 -5.670 41.390 -5.360 ;
        RECT 41.980 -5.670 42.300 -5.360 ;
        RECT 43.610 -5.590 43.900 -5.330 ;
        RECT 43.680 -5.810 43.820 -5.590 ;
        RECT 45.180 -5.670 45.500 -5.360 ;
        RECT 46.820 -5.670 47.140 -5.360 ;
        RECT 47.730 -5.670 48.050 -5.360 ;
        RECT 49.360 -5.590 49.650 -5.330 ;
        RECT 49.430 -5.810 49.570 -5.590 ;
        RECT 50.930 -5.670 51.250 -5.360 ;
        RECT 52.570 -5.670 52.890 -5.360 ;
        RECT 53.480 -5.670 53.800 -5.360 ;
        RECT 55.110 -5.590 55.400 -5.330 ;
        RECT 55.180 -5.810 55.320 -5.590 ;
        RECT 56.680 -5.670 57.000 -5.360 ;
        RECT 58.320 -5.670 58.640 -5.360 ;
        RECT 59.230 -5.670 59.550 -5.360 ;
        RECT 60.860 -5.590 61.150 -5.330 ;
        RECT 60.930 -5.810 61.070 -5.590 ;
        RECT 62.430 -5.670 62.750 -5.360 ;
        RECT 64.070 -5.670 64.390 -5.360 ;
        RECT 64.980 -5.670 65.300 -5.360 ;
        RECT 66.610 -5.590 66.900 -5.330 ;
        RECT 66.680 -5.810 66.820 -5.590 ;
        RECT 68.180 -5.670 68.500 -5.360 ;
        RECT 69.820 -5.670 70.140 -5.360 ;
        RECT 70.730 -5.670 71.050 -5.360 ;
        RECT 72.360 -5.590 72.650 -5.330 ;
        RECT 72.430 -5.810 72.570 -5.590 ;
        RECT 73.930 -5.670 74.250 -5.360 ;
        RECT 75.570 -5.670 75.890 -5.360 ;
        RECT 76.480 -5.670 76.800 -5.360 ;
        RECT 78.110 -5.590 78.400 -5.330 ;
        RECT 78.180 -5.810 78.320 -5.590 ;
        RECT 79.680 -5.670 80.000 -5.360 ;
        RECT 81.320 -5.670 81.640 -5.360 ;
        RECT 82.230 -5.670 82.550 -5.360 ;
        RECT 83.860 -5.590 84.150 -5.330 ;
        RECT 83.930 -5.810 84.070 -5.590 ;
        RECT 85.430 -5.670 85.750 -5.360 ;
        RECT 87.070 -5.670 87.390 -5.360 ;
        RECT 87.980 -5.670 88.300 -5.360 ;
        RECT 89.610 -5.590 89.900 -5.330 ;
        RECT 89.680 -5.810 89.820 -5.590 ;
        RECT 91.180 -5.670 91.500 -5.360 ;
        RECT 92.820 -5.670 93.140 -5.360 ;
        RECT 93.730 -5.670 94.050 -5.360 ;
        RECT 1.260 -5.950 94.660 -5.810 ;
        RECT 1.260 -6.010 1.580 -5.950 ;
        RECT 7.140 -6.240 7.280 -5.950 ;
        RECT 12.890 -6.240 13.030 -5.950 ;
        RECT 18.640 -6.240 18.780 -5.950 ;
        RECT 24.390 -6.240 24.530 -5.950 ;
        RECT 30.140 -6.240 30.280 -5.950 ;
        RECT 35.890 -6.240 36.030 -5.950 ;
        RECT 41.640 -6.240 41.780 -5.950 ;
        RECT 47.390 -6.240 47.530 -5.950 ;
        RECT 53.140 -6.240 53.280 -5.950 ;
        RECT 58.890 -6.240 59.030 -5.950 ;
        RECT 64.640 -6.240 64.780 -5.950 ;
        RECT 70.390 -6.240 70.530 -5.950 ;
        RECT 76.140 -6.240 76.280 -5.950 ;
        RECT 81.890 -6.240 82.030 -5.950 ;
        RECT 87.640 -6.240 87.780 -5.950 ;
        RECT 93.390 -6.240 93.530 -5.950 ;
        RECT 7.060 -6.490 7.350 -6.240 ;
        RECT 12.810 -6.490 13.100 -6.240 ;
        RECT 18.560 -6.490 18.850 -6.240 ;
        RECT 24.310 -6.490 24.600 -6.240 ;
        RECT 30.060 -6.490 30.350 -6.240 ;
        RECT 35.810 -6.490 36.100 -6.240 ;
        RECT 41.560 -6.490 41.850 -6.240 ;
        RECT 47.310 -6.490 47.600 -6.240 ;
        RECT 53.060 -6.490 53.350 -6.240 ;
        RECT 58.810 -6.490 59.100 -6.240 ;
        RECT 64.560 -6.490 64.850 -6.240 ;
        RECT 70.310 -6.490 70.600 -6.240 ;
        RECT 76.060 -6.490 76.350 -6.240 ;
        RECT 81.810 -6.490 82.100 -6.240 ;
        RECT 87.560 -6.490 87.850 -6.240 ;
        RECT 93.310 -6.490 93.600 -6.240 ;
        RECT 2.960 -7.000 3.280 -6.690 ;
        RECT 3.870 -7.000 4.190 -6.690 ;
        RECT 5.460 -7.090 5.830 -6.780 ;
        RECT 8.710 -7.000 9.030 -6.690 ;
        RECT 9.620 -7.000 9.940 -6.690 ;
        RECT 11.210 -7.090 11.580 -6.780 ;
        RECT 14.460 -7.000 14.780 -6.690 ;
        RECT 15.370 -7.000 15.690 -6.690 ;
        RECT 16.960 -7.090 17.330 -6.780 ;
        RECT 20.210 -7.000 20.530 -6.690 ;
        RECT 21.120 -7.000 21.440 -6.690 ;
        RECT 22.710 -7.090 23.080 -6.780 ;
        RECT 25.960 -7.000 26.280 -6.690 ;
        RECT 26.870 -7.000 27.190 -6.690 ;
        RECT 28.460 -7.090 28.830 -6.780 ;
        RECT 31.710 -7.000 32.030 -6.690 ;
        RECT 32.620 -7.000 32.940 -6.690 ;
        RECT 34.210 -7.090 34.580 -6.780 ;
        RECT 37.460 -7.000 37.780 -6.690 ;
        RECT 38.370 -7.000 38.690 -6.690 ;
        RECT 39.960 -7.090 40.330 -6.780 ;
        RECT 43.210 -7.000 43.530 -6.690 ;
        RECT 44.120 -7.000 44.440 -6.690 ;
        RECT 45.710 -7.090 46.080 -6.780 ;
        RECT 48.960 -7.000 49.280 -6.690 ;
        RECT 49.870 -7.000 50.190 -6.690 ;
        RECT 51.460 -7.090 51.830 -6.780 ;
        RECT 54.710 -7.000 55.030 -6.690 ;
        RECT 55.620 -7.000 55.940 -6.690 ;
        RECT 57.210 -7.090 57.580 -6.780 ;
        RECT 60.460 -7.000 60.780 -6.690 ;
        RECT 61.370 -7.000 61.690 -6.690 ;
        RECT 62.960 -7.090 63.330 -6.780 ;
        RECT 66.210 -7.000 66.530 -6.690 ;
        RECT 67.120 -7.000 67.440 -6.690 ;
        RECT 68.710 -7.090 69.080 -6.780 ;
        RECT 71.960 -7.000 72.280 -6.690 ;
        RECT 72.870 -7.000 73.190 -6.690 ;
        RECT 74.460 -7.090 74.830 -6.780 ;
        RECT 77.710 -7.000 78.030 -6.690 ;
        RECT 78.620 -7.000 78.940 -6.690 ;
        RECT 80.210 -7.090 80.580 -6.780 ;
        RECT 83.460 -7.000 83.780 -6.690 ;
        RECT 84.370 -7.000 84.690 -6.690 ;
        RECT 85.960 -7.090 86.330 -6.780 ;
        RECT 89.210 -7.000 89.530 -6.690 ;
        RECT 90.120 -7.000 90.440 -6.690 ;
        RECT 91.710 -7.090 92.080 -6.780 ;
        RECT 1.260 -7.230 1.580 -7.150 ;
        RECT 2.460 -7.230 2.760 -7.170 ;
        RECT 8.210 -7.230 8.510 -7.170 ;
        RECT 13.960 -7.230 14.260 -7.170 ;
        RECT 19.710 -7.230 20.010 -7.170 ;
        RECT 25.460 -7.230 25.760 -7.170 ;
        RECT 31.210 -7.230 31.510 -7.170 ;
        RECT 36.960 -7.230 37.260 -7.170 ;
        RECT 42.710 -7.230 43.010 -7.170 ;
        RECT 48.460 -7.230 48.760 -7.170 ;
        RECT 54.210 -7.230 54.510 -7.170 ;
        RECT 59.960 -7.230 60.260 -7.170 ;
        RECT 65.710 -7.230 66.010 -7.170 ;
        RECT 71.460 -7.230 71.760 -7.170 ;
        RECT 77.210 -7.230 77.510 -7.170 ;
        RECT 82.960 -7.230 83.260 -7.170 ;
        RECT 88.710 -7.230 89.010 -7.170 ;
        RECT 1.260 -7.370 94.660 -7.230 ;
        RECT 1.260 -7.470 1.580 -7.370 ;
        RECT 2.460 -7.450 2.760 -7.370 ;
        RECT 8.210 -7.450 8.510 -7.370 ;
        RECT 13.960 -7.450 14.260 -7.370 ;
        RECT 19.710 -7.450 20.010 -7.370 ;
        RECT 25.460 -7.450 25.760 -7.370 ;
        RECT 31.210 -7.450 31.510 -7.370 ;
        RECT 36.960 -7.450 37.260 -7.370 ;
        RECT 42.710 -7.450 43.010 -7.370 ;
        RECT 48.460 -7.450 48.760 -7.370 ;
        RECT 54.210 -7.450 54.510 -7.370 ;
        RECT 59.960 -7.450 60.260 -7.370 ;
        RECT 65.710 -7.450 66.010 -7.370 ;
        RECT 71.460 -7.450 71.760 -7.370 ;
        RECT 77.210 -7.450 77.510 -7.370 ;
        RECT 82.960 -7.450 83.260 -7.370 ;
        RECT 88.710 -7.450 89.010 -7.370 ;
        RECT 1.260 -8.040 1.580 -7.950 ;
        RECT 8.010 -8.040 8.310 -7.940 ;
        RECT 13.760 -8.040 14.060 -7.940 ;
        RECT 19.510 -8.040 19.810 -7.940 ;
        RECT 25.260 -8.040 25.560 -7.940 ;
        RECT 31.010 -8.040 31.310 -7.940 ;
        RECT 36.760 -8.040 37.060 -7.940 ;
        RECT 42.510 -8.040 42.810 -7.940 ;
        RECT 48.260 -8.040 48.560 -7.940 ;
        RECT 54.010 -8.040 54.310 -7.940 ;
        RECT 59.760 -8.040 60.060 -7.940 ;
        RECT 65.510 -8.040 65.810 -7.940 ;
        RECT 71.260 -8.040 71.560 -7.940 ;
        RECT 77.010 -8.040 77.310 -7.940 ;
        RECT 82.760 -8.040 83.060 -7.940 ;
        RECT 88.510 -8.040 88.810 -7.940 ;
        RECT 94.260 -8.040 94.560 -7.940 ;
        RECT 1.260 -8.180 94.660 -8.040 ;
        RECT 1.260 -8.270 1.580 -8.180 ;
        RECT 8.010 -8.270 8.310 -8.180 ;
        RECT 13.760 -8.270 14.060 -8.180 ;
        RECT 19.510 -8.270 19.810 -8.180 ;
        RECT 25.260 -8.270 25.560 -8.180 ;
        RECT 31.010 -8.270 31.310 -8.180 ;
        RECT 36.760 -8.270 37.060 -8.180 ;
        RECT 42.510 -8.270 42.810 -8.180 ;
        RECT 48.260 -8.270 48.560 -8.180 ;
        RECT 54.010 -8.270 54.310 -8.180 ;
        RECT 59.760 -8.270 60.060 -8.180 ;
        RECT 65.510 -8.270 65.810 -8.180 ;
        RECT 71.260 -8.270 71.560 -8.180 ;
        RECT 77.010 -8.270 77.310 -8.180 ;
        RECT 82.760 -8.270 83.060 -8.180 ;
        RECT 88.510 -8.270 88.810 -8.180 ;
        RECT 94.260 -8.270 94.560 -8.180 ;
        RECT 3.360 -8.590 3.650 -8.330 ;
        RECT 1.260 -8.810 1.580 -8.720 ;
        RECT 3.430 -8.810 3.570 -8.590 ;
        RECT 4.930 -8.670 5.250 -8.360 ;
        RECT 6.570 -8.670 6.890 -8.360 ;
        RECT 7.480 -8.670 7.800 -8.360 ;
        RECT 9.110 -8.590 9.400 -8.330 ;
        RECT 9.180 -8.810 9.320 -8.590 ;
        RECT 10.680 -8.670 11.000 -8.360 ;
        RECT 12.320 -8.670 12.640 -8.360 ;
        RECT 13.230 -8.670 13.550 -8.360 ;
        RECT 14.860 -8.590 15.150 -8.330 ;
        RECT 14.930 -8.810 15.070 -8.590 ;
        RECT 16.430 -8.670 16.750 -8.360 ;
        RECT 18.070 -8.670 18.390 -8.360 ;
        RECT 18.980 -8.670 19.300 -8.360 ;
        RECT 20.610 -8.590 20.900 -8.330 ;
        RECT 20.680 -8.810 20.820 -8.590 ;
        RECT 22.180 -8.670 22.500 -8.360 ;
        RECT 23.820 -8.670 24.140 -8.360 ;
        RECT 24.730 -8.670 25.050 -8.360 ;
        RECT 26.360 -8.590 26.650 -8.330 ;
        RECT 26.430 -8.810 26.570 -8.590 ;
        RECT 27.930 -8.670 28.250 -8.360 ;
        RECT 29.570 -8.670 29.890 -8.360 ;
        RECT 30.480 -8.670 30.800 -8.360 ;
        RECT 32.110 -8.590 32.400 -8.330 ;
        RECT 32.180 -8.810 32.320 -8.590 ;
        RECT 33.680 -8.670 34.000 -8.360 ;
        RECT 35.320 -8.670 35.640 -8.360 ;
        RECT 36.230 -8.670 36.550 -8.360 ;
        RECT 37.860 -8.590 38.150 -8.330 ;
        RECT 37.930 -8.810 38.070 -8.590 ;
        RECT 39.430 -8.670 39.750 -8.360 ;
        RECT 41.070 -8.670 41.390 -8.360 ;
        RECT 41.980 -8.670 42.300 -8.360 ;
        RECT 43.610 -8.590 43.900 -8.330 ;
        RECT 43.680 -8.810 43.820 -8.590 ;
        RECT 45.180 -8.670 45.500 -8.360 ;
        RECT 46.820 -8.670 47.140 -8.360 ;
        RECT 47.730 -8.670 48.050 -8.360 ;
        RECT 49.360 -8.590 49.650 -8.330 ;
        RECT 49.430 -8.810 49.570 -8.590 ;
        RECT 50.930 -8.670 51.250 -8.360 ;
        RECT 52.570 -8.670 52.890 -8.360 ;
        RECT 53.480 -8.670 53.800 -8.360 ;
        RECT 55.110 -8.590 55.400 -8.330 ;
        RECT 55.180 -8.810 55.320 -8.590 ;
        RECT 56.680 -8.670 57.000 -8.360 ;
        RECT 58.320 -8.670 58.640 -8.360 ;
        RECT 59.230 -8.670 59.550 -8.360 ;
        RECT 60.860 -8.590 61.150 -8.330 ;
        RECT 60.930 -8.810 61.070 -8.590 ;
        RECT 62.430 -8.670 62.750 -8.360 ;
        RECT 64.070 -8.670 64.390 -8.360 ;
        RECT 64.980 -8.670 65.300 -8.360 ;
        RECT 66.610 -8.590 66.900 -8.330 ;
        RECT 66.680 -8.810 66.820 -8.590 ;
        RECT 68.180 -8.670 68.500 -8.360 ;
        RECT 69.820 -8.670 70.140 -8.360 ;
        RECT 70.730 -8.670 71.050 -8.360 ;
        RECT 72.360 -8.590 72.650 -8.330 ;
        RECT 72.430 -8.810 72.570 -8.590 ;
        RECT 73.930 -8.670 74.250 -8.360 ;
        RECT 75.570 -8.670 75.890 -8.360 ;
        RECT 76.480 -8.670 76.800 -8.360 ;
        RECT 78.110 -8.590 78.400 -8.330 ;
        RECT 78.180 -8.810 78.320 -8.590 ;
        RECT 79.680 -8.670 80.000 -8.360 ;
        RECT 81.320 -8.670 81.640 -8.360 ;
        RECT 82.230 -8.670 82.550 -8.360 ;
        RECT 83.860 -8.590 84.150 -8.330 ;
        RECT 83.930 -8.810 84.070 -8.590 ;
        RECT 85.430 -8.670 85.750 -8.360 ;
        RECT 87.070 -8.670 87.390 -8.360 ;
        RECT 87.980 -8.670 88.300 -8.360 ;
        RECT 89.610 -8.590 89.900 -8.330 ;
        RECT 89.680 -8.810 89.820 -8.590 ;
        RECT 91.180 -8.670 91.500 -8.360 ;
        RECT 92.820 -8.670 93.140 -8.360 ;
        RECT 93.730 -8.670 94.050 -8.360 ;
        RECT 1.260 -8.950 94.660 -8.810 ;
        RECT 1.260 -9.040 1.580 -8.950 ;
        RECT 2.960 -9.410 3.280 -9.100 ;
        RECT 3.870 -9.410 4.190 -9.100 ;
        RECT 7.060 -9.190 7.350 -8.950 ;
        RECT 5.460 -9.500 5.830 -9.190 ;
        RECT 8.710 -9.410 9.030 -9.100 ;
        RECT 9.620 -9.410 9.940 -9.100 ;
        RECT 12.810 -9.190 13.100 -8.950 ;
        RECT 11.210 -9.500 11.580 -9.190 ;
        RECT 14.460 -9.410 14.780 -9.100 ;
        RECT 15.370 -9.410 15.690 -9.100 ;
        RECT 18.560 -9.190 18.850 -8.950 ;
        RECT 16.960 -9.500 17.330 -9.190 ;
        RECT 20.210 -9.410 20.530 -9.100 ;
        RECT 21.120 -9.410 21.440 -9.100 ;
        RECT 24.310 -9.190 24.600 -8.950 ;
        RECT 22.710 -9.500 23.080 -9.190 ;
        RECT 25.960 -9.410 26.280 -9.100 ;
        RECT 26.870 -9.410 27.190 -9.100 ;
        RECT 30.060 -9.190 30.350 -8.950 ;
        RECT 28.460 -9.500 28.830 -9.190 ;
        RECT 31.710 -9.410 32.030 -9.100 ;
        RECT 32.620 -9.410 32.940 -9.100 ;
        RECT 35.810 -9.190 36.100 -8.950 ;
        RECT 34.210 -9.500 34.580 -9.190 ;
        RECT 37.460 -9.410 37.780 -9.100 ;
        RECT 38.370 -9.410 38.690 -9.100 ;
        RECT 41.560 -9.190 41.850 -8.950 ;
        RECT 39.960 -9.500 40.330 -9.190 ;
        RECT 43.210 -9.410 43.530 -9.100 ;
        RECT 44.120 -9.410 44.440 -9.100 ;
        RECT 47.310 -9.190 47.600 -8.950 ;
        RECT 45.710 -9.500 46.080 -9.190 ;
        RECT 48.960 -9.410 49.280 -9.100 ;
        RECT 49.870 -9.410 50.190 -9.100 ;
        RECT 53.060 -9.190 53.350 -8.950 ;
        RECT 51.460 -9.500 51.830 -9.190 ;
        RECT 54.710 -9.410 55.030 -9.100 ;
        RECT 55.620 -9.410 55.940 -9.100 ;
        RECT 58.810 -9.190 59.100 -8.950 ;
        RECT 57.210 -9.500 57.580 -9.190 ;
        RECT 60.460 -9.410 60.780 -9.100 ;
        RECT 61.370 -9.410 61.690 -9.100 ;
        RECT 64.560 -9.190 64.850 -8.950 ;
        RECT 62.960 -9.500 63.330 -9.190 ;
        RECT 66.210 -9.410 66.530 -9.100 ;
        RECT 67.120 -9.410 67.440 -9.100 ;
        RECT 70.310 -9.190 70.600 -8.950 ;
        RECT 68.710 -9.500 69.080 -9.190 ;
        RECT 71.960 -9.410 72.280 -9.100 ;
        RECT 72.870 -9.410 73.190 -9.100 ;
        RECT 76.060 -9.190 76.350 -8.950 ;
        RECT 74.460 -9.500 74.830 -9.190 ;
        RECT 77.710 -9.410 78.030 -9.100 ;
        RECT 78.620 -9.410 78.940 -9.100 ;
        RECT 81.810 -9.190 82.100 -8.950 ;
        RECT 80.210 -9.500 80.580 -9.190 ;
        RECT 83.460 -9.410 83.780 -9.100 ;
        RECT 84.370 -9.410 84.690 -9.100 ;
        RECT 87.560 -9.190 87.850 -8.950 ;
        RECT 85.960 -9.500 86.330 -9.190 ;
        RECT 89.210 -9.410 89.530 -9.100 ;
        RECT 90.120 -9.410 90.440 -9.100 ;
        RECT 93.310 -9.190 93.600 -8.950 ;
        RECT 91.710 -9.500 92.080 -9.190 ;
        RECT 1.260 -9.640 1.580 -9.520 ;
        RECT 2.460 -9.640 2.760 -9.570 ;
        RECT 8.210 -9.640 8.510 -9.570 ;
        RECT 13.960 -9.640 14.260 -9.570 ;
        RECT 19.710 -9.640 20.010 -9.570 ;
        RECT 25.460 -9.640 25.760 -9.570 ;
        RECT 31.210 -9.640 31.510 -9.570 ;
        RECT 36.960 -9.640 37.260 -9.570 ;
        RECT 42.710 -9.640 43.010 -9.570 ;
        RECT 48.460 -9.640 48.760 -9.570 ;
        RECT 54.210 -9.640 54.510 -9.570 ;
        RECT 59.960 -9.640 60.260 -9.570 ;
        RECT 65.710 -9.640 66.010 -9.570 ;
        RECT 71.460 -9.640 71.760 -9.570 ;
        RECT 77.210 -9.640 77.510 -9.570 ;
        RECT 82.960 -9.640 83.260 -9.570 ;
        RECT 88.710 -9.640 89.010 -9.570 ;
        RECT 1.260 -9.780 94.660 -9.640 ;
        RECT 1.260 -9.840 1.580 -9.780 ;
        RECT 2.460 -9.860 2.760 -9.780 ;
        RECT 8.210 -9.860 8.510 -9.780 ;
        RECT 13.960 -9.860 14.260 -9.780 ;
        RECT 19.710 -9.860 20.010 -9.780 ;
        RECT 25.460 -9.860 25.760 -9.780 ;
        RECT 31.210 -9.860 31.510 -9.780 ;
        RECT 36.960 -9.860 37.260 -9.780 ;
        RECT 42.710 -9.860 43.010 -9.780 ;
        RECT 48.460 -9.860 48.760 -9.780 ;
        RECT 54.210 -9.860 54.510 -9.780 ;
        RECT 59.960 -9.860 60.260 -9.780 ;
        RECT 65.710 -9.860 66.010 -9.780 ;
        RECT 71.460 -9.860 71.760 -9.780 ;
        RECT 77.210 -9.860 77.510 -9.780 ;
        RECT 82.960 -9.860 83.260 -9.780 ;
        RECT 88.710 -9.860 89.010 -9.780 ;
        RECT 1.270 -10.450 1.590 -10.390 ;
        RECT 8.010 -10.450 8.310 -10.350 ;
        RECT 13.760 -10.450 14.060 -10.350 ;
        RECT 19.510 -10.450 19.810 -10.350 ;
        RECT 25.260 -10.450 25.560 -10.350 ;
        RECT 31.010 -10.450 31.310 -10.350 ;
        RECT 36.760 -10.450 37.060 -10.350 ;
        RECT 42.510 -10.450 42.810 -10.350 ;
        RECT 48.260 -10.450 48.560 -10.350 ;
        RECT 54.010 -10.450 54.310 -10.350 ;
        RECT 59.760 -10.450 60.060 -10.350 ;
        RECT 65.510 -10.450 65.810 -10.350 ;
        RECT 71.260 -10.450 71.560 -10.350 ;
        RECT 77.010 -10.450 77.310 -10.350 ;
        RECT 82.760 -10.450 83.060 -10.350 ;
        RECT 88.510 -10.450 88.810 -10.350 ;
        RECT 94.260 -10.450 94.560 -10.350 ;
        RECT 1.270 -10.590 94.660 -10.450 ;
        RECT 1.270 -10.710 1.590 -10.590 ;
        RECT 8.010 -10.680 8.310 -10.590 ;
        RECT 13.760 -10.680 14.060 -10.590 ;
        RECT 19.510 -10.680 19.810 -10.590 ;
        RECT 25.260 -10.680 25.560 -10.590 ;
        RECT 31.010 -10.680 31.310 -10.590 ;
        RECT 36.760 -10.680 37.060 -10.590 ;
        RECT 42.510 -10.680 42.810 -10.590 ;
        RECT 48.260 -10.680 48.560 -10.590 ;
        RECT 54.010 -10.680 54.310 -10.590 ;
        RECT 59.760 -10.680 60.060 -10.590 ;
        RECT 65.510 -10.680 65.810 -10.590 ;
        RECT 71.260 -10.680 71.560 -10.590 ;
        RECT 77.010 -10.680 77.310 -10.590 ;
        RECT 82.760 -10.680 83.060 -10.590 ;
        RECT 88.510 -10.680 88.810 -10.590 ;
        RECT 94.260 -10.680 94.560 -10.590 ;
        RECT 3.360 -11.000 3.650 -10.740 ;
        RECT 1.260 -11.220 1.580 -11.160 ;
        RECT 3.430 -11.220 3.570 -11.000 ;
        RECT 4.930 -11.080 5.250 -10.770 ;
        RECT 6.570 -11.080 6.890 -10.770 ;
        RECT 7.480 -11.080 7.800 -10.770 ;
        RECT 9.110 -11.000 9.400 -10.740 ;
        RECT 9.180 -11.220 9.320 -11.000 ;
        RECT 10.680 -11.080 11.000 -10.770 ;
        RECT 12.320 -11.080 12.640 -10.770 ;
        RECT 13.230 -11.080 13.550 -10.770 ;
        RECT 14.860 -11.000 15.150 -10.740 ;
        RECT 14.930 -11.220 15.070 -11.000 ;
        RECT 16.430 -11.080 16.750 -10.770 ;
        RECT 18.070 -11.080 18.390 -10.770 ;
        RECT 18.980 -11.080 19.300 -10.770 ;
        RECT 20.610 -11.000 20.900 -10.740 ;
        RECT 20.680 -11.220 20.820 -11.000 ;
        RECT 22.180 -11.080 22.500 -10.770 ;
        RECT 23.820 -11.080 24.140 -10.770 ;
        RECT 24.730 -11.080 25.050 -10.770 ;
        RECT 26.360 -11.000 26.650 -10.740 ;
        RECT 26.430 -11.220 26.570 -11.000 ;
        RECT 27.930 -11.080 28.250 -10.770 ;
        RECT 29.570 -11.080 29.890 -10.770 ;
        RECT 30.480 -11.080 30.800 -10.770 ;
        RECT 32.110 -11.000 32.400 -10.740 ;
        RECT 32.180 -11.220 32.320 -11.000 ;
        RECT 33.680 -11.080 34.000 -10.770 ;
        RECT 35.320 -11.080 35.640 -10.770 ;
        RECT 36.230 -11.080 36.550 -10.770 ;
        RECT 37.860 -11.000 38.150 -10.740 ;
        RECT 37.930 -11.220 38.070 -11.000 ;
        RECT 39.430 -11.080 39.750 -10.770 ;
        RECT 41.070 -11.080 41.390 -10.770 ;
        RECT 41.980 -11.080 42.300 -10.770 ;
        RECT 43.610 -11.000 43.900 -10.740 ;
        RECT 43.680 -11.220 43.820 -11.000 ;
        RECT 45.180 -11.080 45.500 -10.770 ;
        RECT 46.820 -11.080 47.140 -10.770 ;
        RECT 47.730 -11.080 48.050 -10.770 ;
        RECT 49.360 -11.000 49.650 -10.740 ;
        RECT 49.430 -11.220 49.570 -11.000 ;
        RECT 50.930 -11.080 51.250 -10.770 ;
        RECT 52.570 -11.080 52.890 -10.770 ;
        RECT 53.480 -11.080 53.800 -10.770 ;
        RECT 55.110 -11.000 55.400 -10.740 ;
        RECT 55.180 -11.220 55.320 -11.000 ;
        RECT 56.680 -11.080 57.000 -10.770 ;
        RECT 58.320 -11.080 58.640 -10.770 ;
        RECT 59.230 -11.080 59.550 -10.770 ;
        RECT 60.860 -11.000 61.150 -10.740 ;
        RECT 60.930 -11.220 61.070 -11.000 ;
        RECT 62.430 -11.080 62.750 -10.770 ;
        RECT 64.070 -11.080 64.390 -10.770 ;
        RECT 64.980 -11.080 65.300 -10.770 ;
        RECT 66.610 -11.000 66.900 -10.740 ;
        RECT 66.680 -11.220 66.820 -11.000 ;
        RECT 68.180 -11.080 68.500 -10.770 ;
        RECT 69.820 -11.080 70.140 -10.770 ;
        RECT 70.730 -11.080 71.050 -10.770 ;
        RECT 72.360 -11.000 72.650 -10.740 ;
        RECT 72.430 -11.220 72.570 -11.000 ;
        RECT 73.930 -11.080 74.250 -10.770 ;
        RECT 75.570 -11.080 75.890 -10.770 ;
        RECT 76.480 -11.080 76.800 -10.770 ;
        RECT 78.110 -11.000 78.400 -10.740 ;
        RECT 78.180 -11.220 78.320 -11.000 ;
        RECT 79.680 -11.080 80.000 -10.770 ;
        RECT 81.320 -11.080 81.640 -10.770 ;
        RECT 82.230 -11.080 82.550 -10.770 ;
        RECT 83.860 -11.000 84.150 -10.740 ;
        RECT 83.930 -11.220 84.070 -11.000 ;
        RECT 85.430 -11.080 85.750 -10.770 ;
        RECT 87.070 -11.080 87.390 -10.770 ;
        RECT 87.980 -11.080 88.300 -10.770 ;
        RECT 89.610 -11.000 89.900 -10.740 ;
        RECT 89.680 -11.220 89.820 -11.000 ;
        RECT 91.180 -11.080 91.500 -10.770 ;
        RECT 92.820 -11.080 93.140 -10.770 ;
        RECT 93.730 -11.080 94.050 -10.770 ;
        RECT 1.260 -11.360 94.660 -11.220 ;
        RECT 1.260 -11.420 1.580 -11.360 ;
        RECT 3.580 -12.680 3.830 -12.560 ;
        RECT 5.230 -12.680 5.550 -12.590 ;
        RECT 6.920 -12.680 7.170 -12.590 ;
        RECT 3.580 -12.820 7.170 -12.680 ;
        RECT 3.580 -12.920 3.830 -12.820 ;
        RECT 5.230 -12.910 5.550 -12.820 ;
        RECT 6.920 -12.910 7.170 -12.820 ;
        RECT 9.330 -12.680 9.580 -12.560 ;
        RECT 10.980 -12.680 11.300 -12.590 ;
        RECT 12.670 -12.680 12.920 -12.590 ;
        RECT 9.330 -12.820 12.920 -12.680 ;
        RECT 9.330 -12.920 9.580 -12.820 ;
        RECT 10.980 -12.910 11.300 -12.820 ;
        RECT 12.670 -12.910 12.920 -12.820 ;
        RECT 15.080 -12.680 15.330 -12.560 ;
        RECT 16.730 -12.680 17.050 -12.590 ;
        RECT 18.420 -12.680 18.670 -12.590 ;
        RECT 15.080 -12.820 18.670 -12.680 ;
        RECT 15.080 -12.920 15.330 -12.820 ;
        RECT 16.730 -12.910 17.050 -12.820 ;
        RECT 18.420 -12.910 18.670 -12.820 ;
        RECT 20.830 -12.680 21.080 -12.560 ;
        RECT 22.480 -12.680 22.800 -12.590 ;
        RECT 24.170 -12.680 24.420 -12.590 ;
        RECT 20.830 -12.820 24.420 -12.680 ;
        RECT 20.830 -12.920 21.080 -12.820 ;
        RECT 22.480 -12.910 22.800 -12.820 ;
        RECT 24.170 -12.910 24.420 -12.820 ;
        RECT 26.580 -12.680 26.830 -12.560 ;
        RECT 28.230 -12.680 28.550 -12.590 ;
        RECT 29.920 -12.680 30.170 -12.590 ;
        RECT 26.580 -12.820 30.170 -12.680 ;
        RECT 26.580 -12.920 26.830 -12.820 ;
        RECT 28.230 -12.910 28.550 -12.820 ;
        RECT 29.920 -12.910 30.170 -12.820 ;
        RECT 32.330 -12.680 32.580 -12.560 ;
        RECT 33.980 -12.680 34.300 -12.590 ;
        RECT 35.670 -12.680 35.920 -12.590 ;
        RECT 32.330 -12.820 35.920 -12.680 ;
        RECT 32.330 -12.920 32.580 -12.820 ;
        RECT 33.980 -12.910 34.300 -12.820 ;
        RECT 35.670 -12.910 35.920 -12.820 ;
        RECT 38.080 -12.680 38.330 -12.560 ;
        RECT 39.730 -12.680 40.050 -12.590 ;
        RECT 41.420 -12.680 41.670 -12.590 ;
        RECT 38.080 -12.820 41.670 -12.680 ;
        RECT 38.080 -12.920 38.330 -12.820 ;
        RECT 39.730 -12.910 40.050 -12.820 ;
        RECT 41.420 -12.910 41.670 -12.820 ;
        RECT 43.830 -12.680 44.080 -12.560 ;
        RECT 45.480 -12.680 45.800 -12.590 ;
        RECT 47.170 -12.680 47.420 -12.590 ;
        RECT 43.830 -12.820 47.420 -12.680 ;
        RECT 43.830 -12.920 44.080 -12.820 ;
        RECT 45.480 -12.910 45.800 -12.820 ;
        RECT 47.170 -12.910 47.420 -12.820 ;
        RECT 49.580 -12.680 49.830 -12.560 ;
        RECT 51.230 -12.680 51.550 -12.590 ;
        RECT 52.920 -12.680 53.170 -12.590 ;
        RECT 49.580 -12.820 53.170 -12.680 ;
        RECT 49.580 -12.920 49.830 -12.820 ;
        RECT 51.230 -12.910 51.550 -12.820 ;
        RECT 52.920 -12.910 53.170 -12.820 ;
        RECT 55.330 -12.680 55.580 -12.560 ;
        RECT 56.980 -12.680 57.300 -12.590 ;
        RECT 58.670 -12.680 58.920 -12.590 ;
        RECT 55.330 -12.820 58.920 -12.680 ;
        RECT 55.330 -12.920 55.580 -12.820 ;
        RECT 56.980 -12.910 57.300 -12.820 ;
        RECT 58.670 -12.910 58.920 -12.820 ;
        RECT 61.080 -12.680 61.330 -12.560 ;
        RECT 62.730 -12.680 63.050 -12.590 ;
        RECT 64.420 -12.680 64.670 -12.590 ;
        RECT 61.080 -12.820 64.670 -12.680 ;
        RECT 61.080 -12.920 61.330 -12.820 ;
        RECT 62.730 -12.910 63.050 -12.820 ;
        RECT 64.420 -12.910 64.670 -12.820 ;
        RECT 66.830 -12.680 67.080 -12.560 ;
        RECT 68.480 -12.680 68.800 -12.590 ;
        RECT 70.170 -12.680 70.420 -12.590 ;
        RECT 66.830 -12.820 70.420 -12.680 ;
        RECT 66.830 -12.920 67.080 -12.820 ;
        RECT 68.480 -12.910 68.800 -12.820 ;
        RECT 70.170 -12.910 70.420 -12.820 ;
        RECT 72.580 -12.680 72.830 -12.560 ;
        RECT 74.230 -12.680 74.550 -12.590 ;
        RECT 75.920 -12.680 76.170 -12.590 ;
        RECT 72.580 -12.820 76.170 -12.680 ;
        RECT 72.580 -12.920 72.830 -12.820 ;
        RECT 74.230 -12.910 74.550 -12.820 ;
        RECT 75.920 -12.910 76.170 -12.820 ;
        RECT 78.330 -12.680 78.580 -12.560 ;
        RECT 79.980 -12.680 80.300 -12.590 ;
        RECT 81.670 -12.680 81.920 -12.590 ;
        RECT 78.330 -12.820 81.920 -12.680 ;
        RECT 78.330 -12.920 78.580 -12.820 ;
        RECT 79.980 -12.910 80.300 -12.820 ;
        RECT 81.670 -12.910 81.920 -12.820 ;
        RECT 84.080 -12.680 84.330 -12.560 ;
        RECT 85.730 -12.680 86.050 -12.590 ;
        RECT 87.420 -12.680 87.670 -12.590 ;
        RECT 84.080 -12.820 87.670 -12.680 ;
        RECT 84.080 -12.920 84.330 -12.820 ;
        RECT 85.730 -12.910 86.050 -12.820 ;
        RECT 87.420 -12.910 87.670 -12.820 ;
        RECT 89.830 -12.680 90.080 -12.560 ;
        RECT 91.480 -12.680 91.800 -12.590 ;
        RECT 93.170 -12.680 93.420 -12.590 ;
        RECT 89.830 -12.820 93.420 -12.680 ;
        RECT 89.830 -12.920 90.080 -12.820 ;
        RECT 91.480 -12.910 91.800 -12.820 ;
        RECT 93.170 -12.910 93.420 -12.820 ;
        RECT 5.940 -14.150 6.260 -13.830 ;
        RECT 11.690 -14.160 12.010 -13.840 ;
        RECT 17.440 -14.180 17.760 -13.860 ;
        RECT 23.190 -14.180 23.510 -13.860 ;
        RECT 28.940 -14.160 29.260 -13.840 ;
        RECT 34.690 -14.130 35.010 -13.810 ;
        RECT 40.400 -14.150 40.800 -13.750 ;
        RECT 46.190 -14.110 46.510 -13.790 ;
        RECT 51.940 -14.160 52.260 -13.840 ;
        RECT 57.690 -14.130 58.010 -13.810 ;
        RECT 63.440 -14.170 63.760 -13.850 ;
        RECT 69.190 -14.180 69.510 -13.860 ;
        RECT 74.940 -14.140 75.260 -13.820 ;
        RECT 80.690 -14.180 81.010 -13.860 ;
        RECT 86.440 -14.140 86.760 -13.820 ;
        RECT 92.190 -14.150 92.510 -13.830 ;
        RECT 3.360 -14.570 3.620 -14.240 ;
        RECT 3.900 -14.570 4.160 -14.240 ;
        RECT 6.610 -14.570 6.870 -14.240 ;
        RECT 7.150 -14.570 7.410 -14.240 ;
        RECT 9.110 -14.570 9.370 -14.240 ;
        RECT 9.650 -14.570 9.910 -14.240 ;
        RECT 12.360 -14.570 12.620 -14.240 ;
        RECT 12.900 -14.570 13.160 -14.240 ;
        RECT 14.860 -14.570 15.120 -14.240 ;
        RECT 15.400 -14.570 15.660 -14.240 ;
        RECT 18.110 -14.570 18.370 -14.240 ;
        RECT 18.650 -14.570 18.910 -14.240 ;
        RECT 20.610 -14.570 20.870 -14.240 ;
        RECT 21.150 -14.570 21.410 -14.240 ;
        RECT 23.860 -14.570 24.120 -14.240 ;
        RECT 24.400 -14.570 24.660 -14.240 ;
        RECT 26.360 -14.570 26.620 -14.240 ;
        RECT 26.900 -14.570 27.160 -14.240 ;
        RECT 29.610 -14.570 29.870 -14.240 ;
        RECT 30.150 -14.570 30.410 -14.240 ;
        RECT 32.110 -14.570 32.370 -14.240 ;
        RECT 32.650 -14.570 32.910 -14.240 ;
        RECT 35.360 -14.570 35.620 -14.240 ;
        RECT 35.900 -14.570 36.160 -14.240 ;
        RECT 37.860 -14.570 38.120 -14.240 ;
        RECT 38.400 -14.570 38.660 -14.240 ;
        RECT 41.110 -14.570 41.370 -14.240 ;
        RECT 41.650 -14.570 41.910 -14.240 ;
        RECT 43.610 -14.570 43.870 -14.240 ;
        RECT 44.150 -14.570 44.410 -14.240 ;
        RECT 46.860 -14.570 47.120 -14.240 ;
        RECT 47.400 -14.570 47.660 -14.240 ;
        RECT 49.360 -14.570 49.620 -14.240 ;
        RECT 49.900 -14.570 50.160 -14.240 ;
        RECT 52.610 -14.570 52.870 -14.240 ;
        RECT 53.150 -14.570 53.410 -14.240 ;
        RECT 55.110 -14.570 55.370 -14.240 ;
        RECT 55.650 -14.570 55.910 -14.240 ;
        RECT 58.360 -14.570 58.620 -14.240 ;
        RECT 58.900 -14.570 59.160 -14.240 ;
        RECT 60.860 -14.570 61.120 -14.240 ;
        RECT 61.400 -14.570 61.660 -14.240 ;
        RECT 64.110 -14.570 64.370 -14.240 ;
        RECT 64.650 -14.570 64.910 -14.240 ;
        RECT 66.610 -14.570 66.870 -14.240 ;
        RECT 67.150 -14.570 67.410 -14.240 ;
        RECT 69.860 -14.570 70.120 -14.240 ;
        RECT 70.400 -14.570 70.660 -14.240 ;
        RECT 72.360 -14.570 72.620 -14.240 ;
        RECT 72.900 -14.570 73.160 -14.240 ;
        RECT 75.610 -14.570 75.870 -14.240 ;
        RECT 76.150 -14.570 76.410 -14.240 ;
        RECT 78.110 -14.570 78.370 -14.240 ;
        RECT 78.650 -14.570 78.910 -14.240 ;
        RECT 81.360 -14.570 81.620 -14.240 ;
        RECT 81.900 -14.570 82.160 -14.240 ;
        RECT 83.860 -14.570 84.120 -14.240 ;
        RECT 84.400 -14.570 84.660 -14.240 ;
        RECT 87.110 -14.570 87.370 -14.240 ;
        RECT 87.650 -14.570 87.910 -14.240 ;
        RECT 89.610 -14.570 89.870 -14.240 ;
        RECT 90.150 -14.570 90.410 -14.240 ;
        RECT 92.860 -14.570 93.120 -14.240 ;
        RECT 93.400 -14.570 93.660 -14.240 ;
        RECT 4.020 -16.040 4.310 -15.990 ;
        RECT 4.980 -16.040 5.270 -15.990 ;
        RECT 4.020 -16.180 5.270 -16.040 ;
        RECT 4.020 -16.240 4.310 -16.180 ;
        RECT 4.980 -16.240 5.270 -16.180 ;
        RECT 9.770 -16.040 10.060 -15.990 ;
        RECT 10.730 -16.040 11.020 -15.990 ;
        RECT 9.770 -16.180 11.020 -16.040 ;
        RECT 9.770 -16.240 10.060 -16.180 ;
        RECT 10.730 -16.240 11.020 -16.180 ;
        RECT 15.520 -16.040 15.810 -15.990 ;
        RECT 16.480 -16.040 16.770 -15.990 ;
        RECT 15.520 -16.180 16.770 -16.040 ;
        RECT 15.520 -16.240 15.810 -16.180 ;
        RECT 16.480 -16.240 16.770 -16.180 ;
        RECT 21.270 -16.040 21.560 -15.990 ;
        RECT 22.230 -16.040 22.520 -15.990 ;
        RECT 21.270 -16.180 22.520 -16.040 ;
        RECT 21.270 -16.240 21.560 -16.180 ;
        RECT 22.230 -16.240 22.520 -16.180 ;
        RECT 27.020 -16.040 27.310 -15.990 ;
        RECT 27.980 -16.040 28.270 -15.990 ;
        RECT 27.020 -16.180 28.270 -16.040 ;
        RECT 27.020 -16.240 27.310 -16.180 ;
        RECT 27.980 -16.240 28.270 -16.180 ;
        RECT 32.770 -16.040 33.060 -15.990 ;
        RECT 33.730 -16.040 34.020 -15.990 ;
        RECT 32.770 -16.180 34.020 -16.040 ;
        RECT 32.770 -16.240 33.060 -16.180 ;
        RECT 33.730 -16.240 34.020 -16.180 ;
        RECT 38.520 -16.040 38.810 -15.990 ;
        RECT 39.480 -16.040 39.770 -15.990 ;
        RECT 38.520 -16.180 39.770 -16.040 ;
        RECT 38.520 -16.240 38.810 -16.180 ;
        RECT 39.480 -16.240 39.770 -16.180 ;
        RECT 44.270 -16.040 44.560 -15.990 ;
        RECT 45.230 -16.040 45.520 -15.990 ;
        RECT 44.270 -16.180 45.520 -16.040 ;
        RECT 44.270 -16.240 44.560 -16.180 ;
        RECT 45.230 -16.240 45.520 -16.180 ;
        RECT 50.020 -16.040 50.310 -15.990 ;
        RECT 50.980 -16.040 51.270 -15.990 ;
        RECT 50.020 -16.180 51.270 -16.040 ;
        RECT 50.020 -16.240 50.310 -16.180 ;
        RECT 50.980 -16.240 51.270 -16.180 ;
        RECT 55.770 -16.040 56.060 -15.990 ;
        RECT 56.730 -16.040 57.020 -15.990 ;
        RECT 55.770 -16.180 57.020 -16.040 ;
        RECT 55.770 -16.240 56.060 -16.180 ;
        RECT 56.730 -16.240 57.020 -16.180 ;
        RECT 61.520 -16.040 61.810 -15.990 ;
        RECT 62.480 -16.040 62.770 -15.990 ;
        RECT 61.520 -16.180 62.770 -16.040 ;
        RECT 61.520 -16.240 61.810 -16.180 ;
        RECT 62.480 -16.240 62.770 -16.180 ;
        RECT 67.270 -16.040 67.560 -15.990 ;
        RECT 68.230 -16.040 68.520 -15.990 ;
        RECT 67.270 -16.180 68.520 -16.040 ;
        RECT 67.270 -16.240 67.560 -16.180 ;
        RECT 68.230 -16.240 68.520 -16.180 ;
        RECT 73.020 -16.040 73.310 -15.990 ;
        RECT 73.980 -16.040 74.270 -15.990 ;
        RECT 73.020 -16.180 74.270 -16.040 ;
        RECT 73.020 -16.240 73.310 -16.180 ;
        RECT 73.980 -16.240 74.270 -16.180 ;
        RECT 78.770 -16.040 79.060 -15.990 ;
        RECT 79.730 -16.040 80.020 -15.990 ;
        RECT 78.770 -16.180 80.020 -16.040 ;
        RECT 78.770 -16.240 79.060 -16.180 ;
        RECT 79.730 -16.240 80.020 -16.180 ;
        RECT 84.520 -16.040 84.810 -15.990 ;
        RECT 85.480 -16.040 85.770 -15.990 ;
        RECT 84.520 -16.180 85.770 -16.040 ;
        RECT 84.520 -16.240 84.810 -16.180 ;
        RECT 85.480 -16.240 85.770 -16.180 ;
        RECT 90.270 -16.040 90.560 -15.990 ;
        RECT 91.230 -16.040 91.520 -15.990 ;
        RECT 90.270 -16.180 91.520 -16.040 ;
        RECT 90.270 -16.240 90.560 -16.180 ;
        RECT 91.230 -16.240 91.520 -16.180 ;
        RECT 5.510 -16.850 5.800 -16.800 ;
        RECT 6.470 -16.850 6.760 -16.810 ;
        RECT 5.510 -16.990 6.760 -16.850 ;
        RECT 5.510 -17.050 5.800 -16.990 ;
        RECT 6.470 -17.060 6.760 -16.990 ;
        RECT 11.260 -16.850 11.550 -16.800 ;
        RECT 12.220 -16.850 12.510 -16.810 ;
        RECT 11.260 -16.990 12.510 -16.850 ;
        RECT 11.260 -17.050 11.550 -16.990 ;
        RECT 12.220 -17.060 12.510 -16.990 ;
        RECT 17.010 -16.850 17.300 -16.800 ;
        RECT 17.970 -16.850 18.260 -16.810 ;
        RECT 17.010 -16.990 18.260 -16.850 ;
        RECT 17.010 -17.050 17.300 -16.990 ;
        RECT 17.970 -17.060 18.260 -16.990 ;
        RECT 22.760 -16.850 23.050 -16.800 ;
        RECT 23.720 -16.850 24.010 -16.810 ;
        RECT 22.760 -16.990 24.010 -16.850 ;
        RECT 22.760 -17.050 23.050 -16.990 ;
        RECT 23.720 -17.060 24.010 -16.990 ;
        RECT 28.510 -16.850 28.800 -16.800 ;
        RECT 29.470 -16.850 29.760 -16.810 ;
        RECT 28.510 -16.990 29.760 -16.850 ;
        RECT 28.510 -17.050 28.800 -16.990 ;
        RECT 29.470 -17.060 29.760 -16.990 ;
        RECT 34.260 -16.850 34.550 -16.800 ;
        RECT 35.220 -16.850 35.510 -16.810 ;
        RECT 34.260 -16.990 35.510 -16.850 ;
        RECT 34.260 -17.050 34.550 -16.990 ;
        RECT 35.220 -17.060 35.510 -16.990 ;
        RECT 40.010 -16.850 40.300 -16.800 ;
        RECT 40.970 -16.850 41.260 -16.810 ;
        RECT 40.010 -16.990 41.260 -16.850 ;
        RECT 40.010 -17.050 40.300 -16.990 ;
        RECT 40.970 -17.060 41.260 -16.990 ;
        RECT 45.760 -16.850 46.050 -16.800 ;
        RECT 46.720 -16.850 47.010 -16.810 ;
        RECT 45.760 -16.990 47.010 -16.850 ;
        RECT 45.760 -17.050 46.050 -16.990 ;
        RECT 46.720 -17.060 47.010 -16.990 ;
        RECT 51.510 -16.850 51.800 -16.800 ;
        RECT 52.470 -16.850 52.760 -16.810 ;
        RECT 51.510 -16.990 52.760 -16.850 ;
        RECT 51.510 -17.050 51.800 -16.990 ;
        RECT 52.470 -17.060 52.760 -16.990 ;
        RECT 57.260 -16.850 57.550 -16.800 ;
        RECT 58.220 -16.850 58.510 -16.810 ;
        RECT 57.260 -16.990 58.510 -16.850 ;
        RECT 57.260 -17.050 57.550 -16.990 ;
        RECT 58.220 -17.060 58.510 -16.990 ;
        RECT 63.010 -16.850 63.300 -16.800 ;
        RECT 63.970 -16.850 64.260 -16.810 ;
        RECT 63.010 -16.990 64.260 -16.850 ;
        RECT 63.010 -17.050 63.300 -16.990 ;
        RECT 63.970 -17.060 64.260 -16.990 ;
        RECT 68.760 -16.850 69.050 -16.800 ;
        RECT 69.720 -16.850 70.010 -16.810 ;
        RECT 68.760 -16.990 70.010 -16.850 ;
        RECT 68.760 -17.050 69.050 -16.990 ;
        RECT 69.720 -17.060 70.010 -16.990 ;
        RECT 74.510 -16.850 74.800 -16.800 ;
        RECT 75.470 -16.850 75.760 -16.810 ;
        RECT 74.510 -16.990 75.760 -16.850 ;
        RECT 74.510 -17.050 74.800 -16.990 ;
        RECT 75.470 -17.060 75.760 -16.990 ;
        RECT 80.260 -16.850 80.550 -16.800 ;
        RECT 81.220 -16.850 81.510 -16.810 ;
        RECT 80.260 -16.990 81.510 -16.850 ;
        RECT 80.260 -17.050 80.550 -16.990 ;
        RECT 81.220 -17.060 81.510 -16.990 ;
        RECT 86.010 -16.850 86.300 -16.800 ;
        RECT 86.970 -16.850 87.260 -16.810 ;
        RECT 86.010 -16.990 87.260 -16.850 ;
        RECT 86.010 -17.050 86.300 -16.990 ;
        RECT 86.970 -17.060 87.260 -16.990 ;
        RECT 91.760 -16.850 92.050 -16.800 ;
        RECT 92.720 -16.850 93.010 -16.810 ;
        RECT 91.760 -16.990 93.010 -16.850 ;
        RECT 91.760 -17.050 92.050 -16.990 ;
        RECT 92.720 -17.060 93.010 -16.990 ;
        RECT 3.400 -18.520 3.730 -18.440 ;
        RECT 7.110 -18.520 7.370 -18.450 ;
        RECT 9.150 -18.520 9.480 -18.440 ;
        RECT 12.860 -18.520 13.120 -18.450 ;
        RECT 14.900 -18.520 15.230 -18.440 ;
        RECT 18.610 -18.520 18.870 -18.450 ;
        RECT 20.650 -18.520 20.980 -18.440 ;
        RECT 24.360 -18.520 24.620 -18.450 ;
        RECT 26.400 -18.520 26.730 -18.440 ;
        RECT 30.110 -18.520 30.370 -18.450 ;
        RECT 32.150 -18.520 32.480 -18.440 ;
        RECT 35.860 -18.520 36.120 -18.450 ;
        RECT 37.900 -18.520 38.230 -18.440 ;
        RECT 41.610 -18.520 41.870 -18.450 ;
        RECT 43.650 -18.520 43.980 -18.440 ;
        RECT 47.360 -18.520 47.620 -18.450 ;
        RECT 49.400 -18.520 49.730 -18.440 ;
        RECT 53.110 -18.520 53.370 -18.450 ;
        RECT 55.150 -18.520 55.480 -18.440 ;
        RECT 58.860 -18.520 59.120 -18.450 ;
        RECT 60.900 -18.520 61.230 -18.440 ;
        RECT 64.610 -18.520 64.870 -18.450 ;
        RECT 66.650 -18.520 66.980 -18.440 ;
        RECT 70.360 -18.520 70.620 -18.450 ;
        RECT 72.400 -18.520 72.730 -18.440 ;
        RECT 76.110 -18.520 76.370 -18.450 ;
        RECT 78.150 -18.520 78.480 -18.440 ;
        RECT 81.860 -18.520 82.120 -18.450 ;
        RECT 83.900 -18.520 84.230 -18.440 ;
        RECT 87.610 -18.520 87.870 -18.450 ;
        RECT 89.650 -18.520 89.980 -18.440 ;
        RECT 93.360 -18.520 93.620 -18.450 ;
        RECT -45.490 -18.660 94.660 -18.520 ;
        RECT 3.400 -18.770 3.730 -18.660 ;
        RECT 7.110 -18.780 7.370 -18.660 ;
        RECT 9.150 -18.770 9.480 -18.660 ;
        RECT 12.860 -18.780 13.120 -18.660 ;
        RECT 14.900 -18.770 15.230 -18.660 ;
        RECT 18.610 -18.780 18.870 -18.660 ;
        RECT 20.650 -18.770 20.980 -18.660 ;
        RECT 24.360 -18.780 24.620 -18.660 ;
        RECT 26.400 -18.770 26.730 -18.660 ;
        RECT 30.110 -18.780 30.370 -18.660 ;
        RECT 32.150 -18.770 32.480 -18.660 ;
        RECT 35.860 -18.780 36.120 -18.660 ;
        RECT 37.900 -18.770 38.230 -18.660 ;
        RECT 41.610 -18.780 41.870 -18.660 ;
        RECT 43.650 -18.770 43.980 -18.660 ;
        RECT 47.360 -18.780 47.620 -18.660 ;
        RECT 49.400 -18.770 49.730 -18.660 ;
        RECT 53.110 -18.780 53.370 -18.660 ;
        RECT 55.150 -18.770 55.480 -18.660 ;
        RECT 58.860 -18.780 59.120 -18.660 ;
        RECT 60.900 -18.770 61.230 -18.660 ;
        RECT 64.610 -18.780 64.870 -18.660 ;
        RECT 66.650 -18.770 66.980 -18.660 ;
        RECT 70.360 -18.780 70.620 -18.660 ;
        RECT 72.400 -18.770 72.730 -18.660 ;
        RECT 76.110 -18.780 76.370 -18.660 ;
        RECT 78.150 -18.770 78.480 -18.660 ;
        RECT 81.860 -18.780 82.120 -18.660 ;
        RECT 83.900 -18.770 84.230 -18.660 ;
        RECT 87.610 -18.780 87.870 -18.660 ;
        RECT 89.650 -18.770 89.980 -18.660 ;
        RECT 93.360 -18.780 93.620 -18.660 ;
        RECT 1.260 -18.990 1.580 -18.930 ;
        RECT 5.330 -18.990 5.620 -18.930 ;
        RECT 8.060 -18.990 8.350 -18.900 ;
        RECT 11.080 -18.990 11.370 -18.930 ;
        RECT 13.810 -18.980 14.100 -18.900 ;
        RECT 13.750 -18.990 14.160 -18.980 ;
        RECT 16.830 -18.990 17.120 -18.930 ;
        RECT 19.560 -18.980 19.850 -18.900 ;
        RECT 19.500 -18.990 19.910 -18.980 ;
        RECT 22.580 -18.990 22.870 -18.930 ;
        RECT 25.310 -18.980 25.600 -18.900 ;
        RECT 25.250 -18.990 25.660 -18.980 ;
        RECT 28.330 -18.990 28.620 -18.930 ;
        RECT 31.060 -18.980 31.350 -18.900 ;
        RECT 31.000 -18.990 31.410 -18.980 ;
        RECT 34.080 -18.990 34.370 -18.930 ;
        RECT 36.810 -18.980 37.100 -18.900 ;
        RECT 36.750 -18.990 37.160 -18.980 ;
        RECT 39.830 -18.990 40.120 -18.930 ;
        RECT 42.560 -18.980 42.850 -18.900 ;
        RECT 42.500 -18.990 42.910 -18.980 ;
        RECT 45.580 -18.990 45.870 -18.930 ;
        RECT 48.310 -18.980 48.600 -18.900 ;
        RECT 48.250 -18.990 48.660 -18.980 ;
        RECT 51.330 -18.990 51.620 -18.930 ;
        RECT 54.060 -18.980 54.350 -18.900 ;
        RECT 54.000 -18.990 54.410 -18.980 ;
        RECT 57.080 -18.990 57.370 -18.930 ;
        RECT 59.810 -18.980 60.100 -18.900 ;
        RECT 59.750 -18.990 60.160 -18.980 ;
        RECT 62.830 -18.990 63.120 -18.930 ;
        RECT 65.560 -18.980 65.850 -18.900 ;
        RECT 65.500 -18.990 65.910 -18.980 ;
        RECT 68.580 -18.990 68.870 -18.930 ;
        RECT 71.310 -18.980 71.600 -18.900 ;
        RECT 71.250 -18.990 71.660 -18.980 ;
        RECT 74.330 -18.990 74.620 -18.930 ;
        RECT 77.060 -18.980 77.350 -18.900 ;
        RECT 77.000 -18.990 77.410 -18.980 ;
        RECT 80.080 -18.990 80.370 -18.930 ;
        RECT 82.810 -18.980 83.100 -18.900 ;
        RECT 82.750 -18.990 83.160 -18.980 ;
        RECT 85.830 -18.990 86.120 -18.930 ;
        RECT 88.560 -18.980 88.850 -18.900 ;
        RECT 88.500 -18.990 88.910 -18.980 ;
        RECT 91.580 -18.990 91.870 -18.930 ;
        RECT 94.170 -18.980 94.460 -18.900 ;
        RECT 94.110 -18.990 94.520 -18.980 ;
        RECT 1.260 -19.130 94.660 -18.990 ;
        RECT 1.260 -19.190 1.580 -19.130 ;
        RECT 5.330 -19.170 5.620 -19.130 ;
        RECT 8.060 -19.190 8.350 -19.130 ;
        RECT 11.080 -19.170 11.370 -19.130 ;
        RECT 13.810 -19.190 14.100 -19.130 ;
        RECT 16.830 -19.170 17.120 -19.130 ;
        RECT 19.560 -19.190 19.850 -19.130 ;
        RECT 22.580 -19.170 22.870 -19.130 ;
        RECT 25.310 -19.190 25.600 -19.130 ;
        RECT 28.330 -19.170 28.620 -19.130 ;
        RECT 31.060 -19.190 31.350 -19.130 ;
        RECT 34.080 -19.170 34.370 -19.130 ;
        RECT 36.810 -19.190 37.100 -19.130 ;
        RECT 39.830 -19.170 40.120 -19.130 ;
        RECT 42.560 -19.190 42.850 -19.130 ;
        RECT 45.580 -19.170 45.870 -19.130 ;
        RECT 48.310 -19.190 48.600 -19.130 ;
        RECT 51.330 -19.170 51.620 -19.130 ;
        RECT 54.060 -19.190 54.350 -19.130 ;
        RECT 57.080 -19.170 57.370 -19.130 ;
        RECT 59.810 -19.190 60.100 -19.130 ;
        RECT 62.830 -19.170 63.120 -19.130 ;
        RECT 65.560 -19.190 65.850 -19.130 ;
        RECT 68.580 -19.170 68.870 -19.130 ;
        RECT 71.310 -19.190 71.600 -19.130 ;
        RECT 74.330 -19.170 74.620 -19.130 ;
        RECT 77.060 -19.190 77.350 -19.130 ;
        RECT 80.080 -19.170 80.370 -19.130 ;
        RECT 82.810 -19.190 83.100 -19.130 ;
        RECT 85.830 -19.170 86.120 -19.130 ;
        RECT 88.560 -19.190 88.850 -19.130 ;
        RECT 91.580 -19.170 91.870 -19.130 ;
        RECT 94.170 -19.190 94.460 -19.130 ;
        RECT 4.100 -20.210 4.380 -19.890 ;
        RECT 6.380 -20.210 6.660 -19.890 ;
        RECT 9.850 -20.210 10.130 -19.890 ;
        RECT 12.130 -20.210 12.410 -19.890 ;
        RECT 15.600 -20.210 15.880 -19.890 ;
        RECT 17.880 -20.210 18.160 -19.890 ;
        RECT 21.350 -20.210 21.630 -19.890 ;
        RECT 23.630 -20.210 23.910 -19.890 ;
        RECT 27.100 -20.210 27.380 -19.890 ;
        RECT 29.380 -20.210 29.660 -19.890 ;
        RECT 32.850 -20.210 33.130 -19.890 ;
        RECT 35.130 -20.210 35.410 -19.890 ;
        RECT 38.600 -20.210 38.880 -19.890 ;
        RECT 40.880 -20.210 41.160 -19.890 ;
        RECT 44.350 -20.210 44.630 -19.890 ;
        RECT 46.630 -20.210 46.910 -19.890 ;
        RECT 50.100 -20.210 50.380 -19.890 ;
        RECT 52.380 -20.210 52.660 -19.890 ;
        RECT 55.850 -20.210 56.130 -19.890 ;
        RECT 58.130 -20.210 58.410 -19.890 ;
        RECT 61.600 -20.210 61.880 -19.890 ;
        RECT 63.880 -20.210 64.160 -19.890 ;
        RECT 67.350 -20.210 67.630 -19.890 ;
        RECT 69.630 -20.210 69.910 -19.890 ;
        RECT 73.100 -20.210 73.380 -19.890 ;
        RECT 75.380 -20.210 75.660 -19.890 ;
        RECT 78.850 -20.210 79.130 -19.890 ;
        RECT 81.130 -20.210 81.410 -19.890 ;
        RECT 84.600 -20.210 84.880 -19.890 ;
        RECT 86.880 -20.210 87.160 -19.890 ;
        RECT 90.350 -20.210 90.630 -19.890 ;
        RECT 92.630 -20.210 92.910 -19.890 ;
        RECT -0.400 -20.380 0.000 -20.250 ;
        RECT 1.260 -20.380 1.590 -20.300 ;
        RECT 3.100 -20.380 3.370 -20.300 ;
        RECT 4.970 -20.380 5.240 -20.310 ;
        RECT 5.510 -20.380 5.780 -20.310 ;
        RECT 7.380 -20.380 7.650 -20.300 ;
        RECT 8.850 -20.380 9.120 -20.300 ;
        RECT 10.720 -20.380 10.990 -20.310 ;
        RECT 11.260 -20.380 11.530 -20.310 ;
        RECT 13.130 -20.380 13.400 -20.300 ;
        RECT 14.600 -20.380 14.870 -20.300 ;
        RECT 16.470 -20.380 16.740 -20.310 ;
        RECT 17.010 -20.380 17.280 -20.310 ;
        RECT 18.880 -20.380 19.150 -20.300 ;
        RECT 20.350 -20.380 20.620 -20.300 ;
        RECT 22.220 -20.380 22.490 -20.310 ;
        RECT 22.760 -20.380 23.030 -20.310 ;
        RECT 24.630 -20.380 24.900 -20.300 ;
        RECT 26.100 -20.380 26.370 -20.300 ;
        RECT 27.970 -20.380 28.240 -20.310 ;
        RECT 28.510 -20.380 28.780 -20.310 ;
        RECT 30.380 -20.380 30.650 -20.300 ;
        RECT 31.850 -20.380 32.120 -20.300 ;
        RECT 33.720 -20.380 33.990 -20.310 ;
        RECT 34.260 -20.380 34.530 -20.310 ;
        RECT 36.130 -20.380 36.400 -20.300 ;
        RECT 37.600 -20.380 37.870 -20.300 ;
        RECT 39.470 -20.380 39.740 -20.310 ;
        RECT 40.010 -20.380 40.280 -20.310 ;
        RECT 41.880 -20.380 42.150 -20.300 ;
        RECT 43.350 -20.380 43.620 -20.300 ;
        RECT 45.220 -20.380 45.490 -20.310 ;
        RECT 45.760 -20.380 46.030 -20.310 ;
        RECT 47.630 -20.380 47.900 -20.300 ;
        RECT 49.100 -20.380 49.370 -20.300 ;
        RECT 50.970 -20.380 51.240 -20.310 ;
        RECT 51.510 -20.380 51.780 -20.310 ;
        RECT 53.380 -20.380 53.650 -20.300 ;
        RECT 54.850 -20.380 55.120 -20.300 ;
        RECT 56.720 -20.380 56.990 -20.310 ;
        RECT 57.260 -20.380 57.530 -20.310 ;
        RECT 59.130 -20.380 59.400 -20.300 ;
        RECT 60.600 -20.380 60.870 -20.300 ;
        RECT 62.470 -20.380 62.740 -20.310 ;
        RECT 63.010 -20.380 63.280 -20.310 ;
        RECT 64.880 -20.380 65.150 -20.300 ;
        RECT 66.350 -20.380 66.620 -20.300 ;
        RECT 68.220 -20.380 68.490 -20.310 ;
        RECT 68.760 -20.380 69.030 -20.310 ;
        RECT 70.630 -20.380 70.900 -20.300 ;
        RECT 72.100 -20.380 72.370 -20.300 ;
        RECT 73.970 -20.380 74.240 -20.310 ;
        RECT 74.510 -20.380 74.780 -20.310 ;
        RECT 76.380 -20.380 76.650 -20.300 ;
        RECT 77.850 -20.380 78.120 -20.300 ;
        RECT 79.720 -20.380 79.990 -20.310 ;
        RECT 80.260 -20.380 80.530 -20.310 ;
        RECT 82.130 -20.380 82.400 -20.300 ;
        RECT 83.600 -20.380 83.870 -20.300 ;
        RECT 85.470 -20.380 85.740 -20.310 ;
        RECT 86.010 -20.380 86.280 -20.310 ;
        RECT 87.880 -20.380 88.150 -20.300 ;
        RECT 89.350 -20.380 89.620 -20.300 ;
        RECT 91.220 -20.380 91.490 -20.310 ;
        RECT 91.760 -20.380 92.030 -20.310 ;
        RECT 93.630 -20.380 93.900 -20.300 ;
        RECT -0.400 -20.520 94.660 -20.380 ;
        RECT -0.400 -20.530 1.590 -20.520 ;
        RECT -0.400 -20.650 0.000 -20.530 ;
        RECT 1.260 -20.620 1.590 -20.530 ;
        RECT 3.100 -20.590 3.370 -20.520 ;
        RECT 4.970 -20.600 5.240 -20.520 ;
        RECT 5.510 -20.600 5.780 -20.520 ;
        RECT 7.380 -20.590 7.650 -20.520 ;
        RECT 8.850 -20.590 9.120 -20.520 ;
        RECT 10.720 -20.600 10.990 -20.520 ;
        RECT 11.260 -20.600 11.530 -20.520 ;
        RECT 13.130 -20.590 13.400 -20.520 ;
        RECT 14.600 -20.590 14.870 -20.520 ;
        RECT 16.470 -20.600 16.740 -20.520 ;
        RECT 17.010 -20.600 17.280 -20.520 ;
        RECT 18.880 -20.590 19.150 -20.520 ;
        RECT 20.350 -20.590 20.620 -20.520 ;
        RECT 22.220 -20.600 22.490 -20.520 ;
        RECT 22.760 -20.600 23.030 -20.520 ;
        RECT 24.630 -20.590 24.900 -20.520 ;
        RECT 26.100 -20.590 26.370 -20.520 ;
        RECT 27.970 -20.600 28.240 -20.520 ;
        RECT 28.510 -20.600 28.780 -20.520 ;
        RECT 30.380 -20.590 30.650 -20.520 ;
        RECT 31.850 -20.590 32.120 -20.520 ;
        RECT 33.720 -20.600 33.990 -20.520 ;
        RECT 34.260 -20.600 34.530 -20.520 ;
        RECT 36.130 -20.590 36.400 -20.520 ;
        RECT 37.600 -20.590 37.870 -20.520 ;
        RECT 39.470 -20.600 39.740 -20.520 ;
        RECT 40.010 -20.600 40.280 -20.520 ;
        RECT 41.880 -20.590 42.150 -20.520 ;
        RECT 43.350 -20.590 43.620 -20.520 ;
        RECT 45.220 -20.600 45.490 -20.520 ;
        RECT 45.760 -20.600 46.030 -20.520 ;
        RECT 47.630 -20.590 47.900 -20.520 ;
        RECT 49.100 -20.590 49.370 -20.520 ;
        RECT 50.970 -20.600 51.240 -20.520 ;
        RECT 51.510 -20.600 51.780 -20.520 ;
        RECT 53.380 -20.590 53.650 -20.520 ;
        RECT 54.850 -20.590 55.120 -20.520 ;
        RECT 56.720 -20.600 56.990 -20.520 ;
        RECT 57.260 -20.600 57.530 -20.520 ;
        RECT 59.130 -20.590 59.400 -20.520 ;
        RECT 60.600 -20.590 60.870 -20.520 ;
        RECT 62.470 -20.600 62.740 -20.520 ;
        RECT 63.010 -20.600 63.280 -20.520 ;
        RECT 64.880 -20.590 65.150 -20.520 ;
        RECT 66.350 -20.590 66.620 -20.520 ;
        RECT 68.220 -20.600 68.490 -20.520 ;
        RECT 68.760 -20.600 69.030 -20.520 ;
        RECT 70.630 -20.590 70.900 -20.520 ;
        RECT 72.100 -20.590 72.370 -20.520 ;
        RECT 73.970 -20.600 74.240 -20.520 ;
        RECT 74.510 -20.600 74.780 -20.520 ;
        RECT 76.380 -20.590 76.650 -20.520 ;
        RECT 77.850 -20.590 78.120 -20.520 ;
        RECT 79.720 -20.600 79.990 -20.520 ;
        RECT 80.260 -20.600 80.530 -20.520 ;
        RECT 82.130 -20.590 82.400 -20.520 ;
        RECT 83.600 -20.590 83.870 -20.520 ;
        RECT 85.470 -20.600 85.740 -20.520 ;
        RECT 86.010 -20.600 86.280 -20.520 ;
        RECT 87.880 -20.590 88.150 -20.520 ;
        RECT 89.350 -20.590 89.620 -20.520 ;
        RECT 91.220 -20.600 91.490 -20.520 ;
        RECT 91.760 -20.600 92.030 -20.520 ;
        RECT 93.630 -20.590 93.900 -20.520 ;
        RECT 2.250 -21.070 2.570 -20.980 ;
        RECT 3.040 -21.070 3.370 -21.010 ;
        RECT 2.250 -21.210 3.370 -21.070 ;
        RECT 2.250 -21.300 2.570 -21.210 ;
        RECT 3.040 -21.260 3.370 -21.210 ;
        RECT 3.580 -21.090 3.870 -21.030 ;
        RECT 5.670 -21.090 6.000 -21.040 ;
        RECT 7.370 -21.090 7.700 -21.030 ;
        RECT 8.060 -21.070 8.380 -20.960 ;
        RECT 8.790 -21.070 9.120 -21.010 ;
        RECT 3.580 -21.230 7.700 -21.090 ;
        RECT 8.000 -21.210 9.120 -21.070 ;
        RECT 3.580 -21.280 3.870 -21.230 ;
        RECT 5.670 -21.280 6.000 -21.230 ;
        RECT 7.370 -21.280 7.700 -21.230 ;
        RECT 8.060 -21.280 8.380 -21.210 ;
        RECT 8.790 -21.260 9.120 -21.210 ;
        RECT 9.330 -21.090 9.620 -21.030 ;
        RECT 11.420 -21.090 11.750 -21.040 ;
        RECT 13.120 -21.090 13.450 -21.030 ;
        RECT 13.780 -21.070 14.100 -20.970 ;
        RECT 14.540 -21.070 14.870 -21.010 ;
        RECT 9.330 -21.230 13.450 -21.090 ;
        RECT 13.750 -21.210 14.870 -21.070 ;
        RECT 9.330 -21.280 9.620 -21.230 ;
        RECT 11.420 -21.280 11.750 -21.230 ;
        RECT 13.120 -21.280 13.450 -21.230 ;
        RECT 13.780 -21.290 14.100 -21.210 ;
        RECT 14.540 -21.260 14.870 -21.210 ;
        RECT 15.080 -21.090 15.370 -21.030 ;
        RECT 17.170 -21.090 17.500 -21.040 ;
        RECT 18.870 -21.090 19.200 -21.030 ;
        RECT 19.560 -21.070 19.880 -20.990 ;
        RECT 20.290 -21.070 20.620 -21.010 ;
        RECT 15.080 -21.230 19.200 -21.090 ;
        RECT 19.500 -21.210 20.620 -21.070 ;
        RECT 15.080 -21.280 15.370 -21.230 ;
        RECT 17.170 -21.280 17.500 -21.230 ;
        RECT 18.870 -21.280 19.200 -21.230 ;
        RECT 19.560 -21.310 19.880 -21.210 ;
        RECT 20.290 -21.260 20.620 -21.210 ;
        RECT 20.830 -21.090 21.120 -21.030 ;
        RECT 22.920 -21.090 23.250 -21.040 ;
        RECT 24.620 -21.090 24.950 -21.030 ;
        RECT 25.310 -21.070 25.630 -20.990 ;
        RECT 26.040 -21.070 26.370 -21.010 ;
        RECT 20.830 -21.230 24.950 -21.090 ;
        RECT 25.250 -21.210 26.370 -21.070 ;
        RECT 20.830 -21.280 21.120 -21.230 ;
        RECT 22.920 -21.280 23.250 -21.230 ;
        RECT 24.620 -21.280 24.950 -21.230 ;
        RECT 25.310 -21.310 25.630 -21.210 ;
        RECT 26.040 -21.260 26.370 -21.210 ;
        RECT 26.580 -21.090 26.870 -21.030 ;
        RECT 28.670 -21.090 29.000 -21.040 ;
        RECT 30.370 -21.090 30.700 -21.030 ;
        RECT 31.020 -21.070 31.340 -21.010 ;
        RECT 31.790 -21.070 32.120 -21.010 ;
        RECT 26.580 -21.230 30.700 -21.090 ;
        RECT 31.000 -21.210 32.120 -21.070 ;
        RECT 26.580 -21.280 26.870 -21.230 ;
        RECT 28.670 -21.280 29.000 -21.230 ;
        RECT 30.370 -21.280 30.700 -21.230 ;
        RECT 31.020 -21.330 31.340 -21.210 ;
        RECT 31.790 -21.260 32.120 -21.210 ;
        RECT 32.330 -21.090 32.620 -21.030 ;
        RECT 34.420 -21.090 34.750 -21.040 ;
        RECT 36.120 -21.090 36.450 -21.030 ;
        RECT 36.790 -21.070 37.110 -21.000 ;
        RECT 37.540 -21.070 37.870 -21.010 ;
        RECT 32.330 -21.230 36.450 -21.090 ;
        RECT 36.750 -21.210 37.870 -21.070 ;
        RECT 32.330 -21.280 32.620 -21.230 ;
        RECT 34.420 -21.280 34.750 -21.230 ;
        RECT 36.120 -21.280 36.450 -21.230 ;
        RECT 36.790 -21.320 37.110 -21.210 ;
        RECT 37.540 -21.260 37.870 -21.210 ;
        RECT 38.080 -21.090 38.370 -21.030 ;
        RECT 40.170 -21.090 40.500 -21.040 ;
        RECT 41.870 -21.090 42.200 -21.030 ;
        RECT 42.590 -21.070 42.910 -20.990 ;
        RECT 43.290 -21.070 43.620 -21.010 ;
        RECT 38.080 -21.230 42.200 -21.090 ;
        RECT 42.500 -21.210 43.620 -21.070 ;
        RECT 38.080 -21.280 38.370 -21.230 ;
        RECT 40.170 -21.280 40.500 -21.230 ;
        RECT 41.870 -21.280 42.200 -21.230 ;
        RECT 42.590 -21.310 42.910 -21.210 ;
        RECT 43.290 -21.260 43.620 -21.210 ;
        RECT 43.830 -21.090 44.120 -21.030 ;
        RECT 45.920 -21.090 46.250 -21.040 ;
        RECT 47.620 -21.090 47.950 -21.030 ;
        RECT 48.290 -21.070 48.610 -20.980 ;
        RECT 49.040 -21.070 49.370 -21.010 ;
        RECT 43.830 -21.230 47.950 -21.090 ;
        RECT 48.250 -21.210 49.370 -21.070 ;
        RECT 43.830 -21.280 44.120 -21.230 ;
        RECT 45.920 -21.280 46.250 -21.230 ;
        RECT 47.620 -21.280 47.950 -21.230 ;
        RECT 48.290 -21.300 48.610 -21.210 ;
        RECT 49.040 -21.260 49.370 -21.210 ;
        RECT 49.580 -21.090 49.870 -21.030 ;
        RECT 51.670 -21.090 52.000 -21.040 ;
        RECT 53.370 -21.090 53.700 -21.030 ;
        RECT 54.060 -21.070 54.380 -21.000 ;
        RECT 54.790 -21.070 55.120 -21.010 ;
        RECT 49.580 -21.230 53.700 -21.090 ;
        RECT 54.000 -21.210 55.120 -21.070 ;
        RECT 49.580 -21.280 49.870 -21.230 ;
        RECT 51.670 -21.280 52.000 -21.230 ;
        RECT 53.370 -21.280 53.700 -21.230 ;
        RECT 54.060 -21.320 54.380 -21.210 ;
        RECT 54.790 -21.260 55.120 -21.210 ;
        RECT 55.330 -21.090 55.620 -21.030 ;
        RECT 57.420 -21.090 57.750 -21.040 ;
        RECT 59.120 -21.090 59.450 -21.030 ;
        RECT 59.800 -21.070 60.120 -20.980 ;
        RECT 60.540 -21.070 60.870 -21.010 ;
        RECT 55.330 -21.230 59.450 -21.090 ;
        RECT 59.750 -21.210 60.870 -21.070 ;
        RECT 55.330 -21.280 55.620 -21.230 ;
        RECT 57.420 -21.280 57.750 -21.230 ;
        RECT 59.120 -21.280 59.450 -21.230 ;
        RECT 59.800 -21.300 60.120 -21.210 ;
        RECT 60.540 -21.260 60.870 -21.210 ;
        RECT 61.080 -21.090 61.370 -21.030 ;
        RECT 63.170 -21.090 63.500 -21.040 ;
        RECT 64.870 -21.090 65.200 -21.030 ;
        RECT 65.530 -21.070 65.850 -20.990 ;
        RECT 66.290 -21.070 66.620 -21.010 ;
        RECT 61.080 -21.230 65.200 -21.090 ;
        RECT 65.500 -21.210 66.620 -21.070 ;
        RECT 61.080 -21.280 61.370 -21.230 ;
        RECT 63.170 -21.280 63.500 -21.230 ;
        RECT 64.870 -21.280 65.200 -21.230 ;
        RECT 65.530 -21.310 65.850 -21.210 ;
        RECT 66.290 -21.260 66.620 -21.210 ;
        RECT 66.830 -21.090 67.120 -21.030 ;
        RECT 68.920 -21.090 69.250 -21.040 ;
        RECT 70.620 -21.090 70.950 -21.030 ;
        RECT 71.300 -21.070 71.620 -21.000 ;
        RECT 72.040 -21.070 72.370 -21.010 ;
        RECT 66.830 -21.230 70.950 -21.090 ;
        RECT 71.250 -21.210 72.370 -21.070 ;
        RECT 66.830 -21.280 67.120 -21.230 ;
        RECT 68.920 -21.280 69.250 -21.230 ;
        RECT 70.620 -21.280 70.950 -21.230 ;
        RECT 71.300 -21.320 71.620 -21.210 ;
        RECT 72.040 -21.260 72.370 -21.210 ;
        RECT 72.580 -21.090 72.870 -21.030 ;
        RECT 74.670 -21.090 75.000 -21.040 ;
        RECT 76.370 -21.090 76.700 -21.030 ;
        RECT 77.060 -21.070 77.380 -21.000 ;
        RECT 77.790 -21.070 78.120 -21.010 ;
        RECT 72.580 -21.230 76.700 -21.090 ;
        RECT 77.000 -21.210 78.120 -21.070 ;
        RECT 72.580 -21.280 72.870 -21.230 ;
        RECT 74.670 -21.280 75.000 -21.230 ;
        RECT 76.370 -21.280 76.700 -21.230 ;
        RECT 77.060 -21.320 77.380 -21.210 ;
        RECT 77.790 -21.260 78.120 -21.210 ;
        RECT 78.330 -21.090 78.620 -21.030 ;
        RECT 80.420 -21.090 80.750 -21.040 ;
        RECT 82.120 -21.090 82.450 -21.030 ;
        RECT 82.790 -21.070 83.110 -21.020 ;
        RECT 83.540 -21.070 83.870 -21.010 ;
        RECT 78.330 -21.230 82.450 -21.090 ;
        RECT 82.750 -21.210 83.870 -21.070 ;
        RECT 78.330 -21.280 78.620 -21.230 ;
        RECT 80.420 -21.280 80.750 -21.230 ;
        RECT 82.120 -21.280 82.450 -21.230 ;
        RECT 82.790 -21.340 83.110 -21.210 ;
        RECT 83.540 -21.260 83.870 -21.210 ;
        RECT 84.080 -21.090 84.370 -21.030 ;
        RECT 86.170 -21.090 86.500 -21.040 ;
        RECT 87.870 -21.090 88.200 -21.030 ;
        RECT 88.540 -21.070 88.860 -21.020 ;
        RECT 89.290 -21.070 89.620 -21.010 ;
        RECT 84.080 -21.230 88.200 -21.090 ;
        RECT 88.500 -21.210 89.620 -21.070 ;
        RECT 84.080 -21.280 84.370 -21.230 ;
        RECT 86.170 -21.280 86.500 -21.230 ;
        RECT 87.870 -21.280 88.200 -21.230 ;
        RECT 88.540 -21.340 88.860 -21.210 ;
        RECT 89.290 -21.260 89.620 -21.210 ;
        RECT 89.830 -21.090 90.120 -21.030 ;
        RECT 91.920 -21.090 92.250 -21.040 ;
        RECT 93.620 -21.090 93.950 -21.030 ;
        RECT 89.830 -21.230 93.950 -21.090 ;
        RECT 89.830 -21.280 90.120 -21.230 ;
        RECT 91.920 -21.280 92.250 -21.230 ;
        RECT 93.620 -21.280 93.950 -21.230 ;
        RECT 3.100 -21.870 3.370 -21.780 ;
        RECT 5.230 -21.870 5.550 -21.780 ;
        RECT 7.380 -21.870 7.650 -21.780 ;
        RECT 3.100 -22.010 7.650 -21.870 ;
        RECT 3.100 -22.070 3.370 -22.010 ;
        RECT 5.230 -22.100 5.550 -22.010 ;
        RECT 7.380 -22.070 7.650 -22.010 ;
        RECT 8.850 -21.870 9.120 -21.780 ;
        RECT 10.980 -21.870 11.300 -21.780 ;
        RECT 13.130 -21.870 13.400 -21.780 ;
        RECT 8.850 -22.010 13.400 -21.870 ;
        RECT 8.850 -22.070 9.120 -22.010 ;
        RECT 10.980 -22.100 11.300 -22.010 ;
        RECT 13.130 -22.070 13.400 -22.010 ;
        RECT 14.600 -21.870 14.870 -21.780 ;
        RECT 16.730 -21.870 17.050 -21.780 ;
        RECT 18.880 -21.870 19.150 -21.780 ;
        RECT 14.600 -22.010 19.150 -21.870 ;
        RECT 14.600 -22.070 14.870 -22.010 ;
        RECT 16.730 -22.100 17.050 -22.010 ;
        RECT 18.880 -22.070 19.150 -22.010 ;
        RECT 20.350 -21.870 20.620 -21.780 ;
        RECT 22.480 -21.870 22.800 -21.780 ;
        RECT 24.630 -21.870 24.900 -21.780 ;
        RECT 20.350 -22.010 24.900 -21.870 ;
        RECT 20.350 -22.070 20.620 -22.010 ;
        RECT 22.480 -22.100 22.800 -22.010 ;
        RECT 24.630 -22.070 24.900 -22.010 ;
        RECT 26.100 -21.870 26.370 -21.780 ;
        RECT 28.230 -21.870 28.550 -21.780 ;
        RECT 30.380 -21.870 30.650 -21.780 ;
        RECT 26.100 -22.010 30.650 -21.870 ;
        RECT 26.100 -22.070 26.370 -22.010 ;
        RECT 28.230 -22.100 28.550 -22.010 ;
        RECT 30.380 -22.070 30.650 -22.010 ;
        RECT 31.850 -21.870 32.120 -21.780 ;
        RECT 33.980 -21.870 34.300 -21.780 ;
        RECT 36.130 -21.870 36.400 -21.780 ;
        RECT 31.850 -22.010 36.400 -21.870 ;
        RECT 31.850 -22.070 32.120 -22.010 ;
        RECT 33.980 -22.100 34.300 -22.010 ;
        RECT 36.130 -22.070 36.400 -22.010 ;
        RECT 37.600 -21.870 37.870 -21.780 ;
        RECT 39.730 -21.870 40.050 -21.780 ;
        RECT 41.880 -21.870 42.150 -21.780 ;
        RECT 37.600 -22.010 42.150 -21.870 ;
        RECT 37.600 -22.070 37.870 -22.010 ;
        RECT 39.730 -22.100 40.050 -22.010 ;
        RECT 41.880 -22.070 42.150 -22.010 ;
        RECT 43.350 -21.870 43.620 -21.780 ;
        RECT 45.480 -21.870 45.800 -21.780 ;
        RECT 47.630 -21.870 47.900 -21.780 ;
        RECT 43.350 -22.010 47.900 -21.870 ;
        RECT 43.350 -22.070 43.620 -22.010 ;
        RECT 45.480 -22.100 45.800 -22.010 ;
        RECT 47.630 -22.070 47.900 -22.010 ;
        RECT 49.100 -21.870 49.370 -21.780 ;
        RECT 51.230 -21.870 51.550 -21.780 ;
        RECT 53.380 -21.870 53.650 -21.780 ;
        RECT 49.100 -22.010 53.650 -21.870 ;
        RECT 49.100 -22.070 49.370 -22.010 ;
        RECT 51.230 -22.100 51.550 -22.010 ;
        RECT 53.380 -22.070 53.650 -22.010 ;
        RECT 54.850 -21.870 55.120 -21.780 ;
        RECT 56.980 -21.870 57.300 -21.780 ;
        RECT 59.130 -21.870 59.400 -21.780 ;
        RECT 54.850 -22.010 59.400 -21.870 ;
        RECT 54.850 -22.070 55.120 -22.010 ;
        RECT 56.980 -22.100 57.300 -22.010 ;
        RECT 59.130 -22.070 59.400 -22.010 ;
        RECT 60.600 -21.870 60.870 -21.780 ;
        RECT 62.730 -21.870 63.050 -21.780 ;
        RECT 64.880 -21.870 65.150 -21.780 ;
        RECT 60.600 -22.010 65.150 -21.870 ;
        RECT 60.600 -22.070 60.870 -22.010 ;
        RECT 62.730 -22.100 63.050 -22.010 ;
        RECT 64.880 -22.070 65.150 -22.010 ;
        RECT 66.350 -21.870 66.620 -21.780 ;
        RECT 68.480 -21.870 68.800 -21.780 ;
        RECT 70.630 -21.870 70.900 -21.780 ;
        RECT 66.350 -22.010 70.900 -21.870 ;
        RECT 66.350 -22.070 66.620 -22.010 ;
        RECT 68.480 -22.100 68.800 -22.010 ;
        RECT 70.630 -22.070 70.900 -22.010 ;
        RECT 72.100 -21.870 72.370 -21.780 ;
        RECT 74.230 -21.870 74.550 -21.780 ;
        RECT 76.380 -21.870 76.650 -21.780 ;
        RECT 72.100 -22.010 76.650 -21.870 ;
        RECT 72.100 -22.070 72.370 -22.010 ;
        RECT 74.230 -22.100 74.550 -22.010 ;
        RECT 76.380 -22.070 76.650 -22.010 ;
        RECT 77.850 -21.870 78.120 -21.780 ;
        RECT 79.980 -21.870 80.300 -21.780 ;
        RECT 82.130 -21.870 82.400 -21.780 ;
        RECT 77.850 -22.010 82.400 -21.870 ;
        RECT 77.850 -22.070 78.120 -22.010 ;
        RECT 79.980 -22.100 80.300 -22.010 ;
        RECT 82.130 -22.070 82.400 -22.010 ;
        RECT 83.600 -21.870 83.870 -21.780 ;
        RECT 85.730 -21.870 86.050 -21.780 ;
        RECT 87.880 -21.870 88.150 -21.780 ;
        RECT 83.600 -22.010 88.150 -21.870 ;
        RECT 83.600 -22.070 83.870 -22.010 ;
        RECT 85.730 -22.100 86.050 -22.010 ;
        RECT 87.880 -22.070 88.150 -22.010 ;
        RECT 89.350 -21.870 89.620 -21.780 ;
        RECT 91.480 -21.870 91.800 -21.780 ;
        RECT 93.630 -21.870 93.900 -21.780 ;
        RECT 89.350 -22.010 93.900 -21.870 ;
        RECT 89.350 -22.070 89.620 -22.010 ;
        RECT 91.480 -22.100 91.800 -22.010 ;
        RECT 93.630 -22.070 93.900 -22.010 ;
        RECT 2.960 -22.800 3.280 -22.740 ;
        RECT 6.620 -22.800 6.910 -22.770 ;
        RECT 7.490 -22.800 7.810 -22.740 ;
        RECT 2.960 -22.940 7.810 -22.800 ;
        RECT 2.960 -23.000 3.280 -22.940 ;
        RECT 6.620 -23.000 6.910 -22.940 ;
        RECT 7.490 -23.000 7.810 -22.940 ;
        RECT 8.710 -22.800 9.030 -22.740 ;
        RECT 9.610 -22.800 9.900 -22.770 ;
        RECT 13.240 -22.800 13.560 -22.740 ;
        RECT 8.710 -22.940 13.560 -22.800 ;
        RECT 8.710 -23.000 9.030 -22.940 ;
        RECT 9.610 -23.000 9.900 -22.940 ;
        RECT 13.240 -23.000 13.560 -22.940 ;
        RECT 14.460 -22.800 14.780 -22.740 ;
        RECT 18.130 -22.800 18.420 -22.770 ;
        RECT 18.990 -22.800 19.310 -22.740 ;
        RECT 14.460 -22.940 19.310 -22.800 ;
        RECT 14.460 -23.000 14.780 -22.940 ;
        RECT 18.130 -23.000 18.420 -22.940 ;
        RECT 18.990 -23.000 19.310 -22.940 ;
        RECT 20.210 -22.800 20.530 -22.740 ;
        RECT 21.110 -22.800 21.400 -22.770 ;
        RECT 24.740 -22.800 25.060 -22.740 ;
        RECT 20.210 -22.940 25.060 -22.800 ;
        RECT 20.210 -23.000 20.530 -22.940 ;
        RECT 21.110 -23.000 21.400 -22.940 ;
        RECT 24.740 -23.000 25.060 -22.940 ;
        RECT 25.960 -22.800 26.280 -22.740 ;
        RECT 29.630 -22.800 29.920 -22.770 ;
        RECT 30.490 -22.800 30.810 -22.740 ;
        RECT 25.960 -22.940 30.810 -22.800 ;
        RECT 25.960 -23.000 26.280 -22.940 ;
        RECT 29.630 -23.000 29.920 -22.940 ;
        RECT 30.490 -23.000 30.810 -22.940 ;
        RECT 31.710 -22.800 32.030 -22.740 ;
        RECT 32.610 -22.800 32.900 -22.770 ;
        RECT 36.240 -22.800 36.560 -22.740 ;
        RECT 31.710 -22.940 36.560 -22.800 ;
        RECT 31.710 -23.000 32.030 -22.940 ;
        RECT 32.610 -23.000 32.900 -22.940 ;
        RECT 36.240 -23.000 36.560 -22.940 ;
        RECT 37.460 -22.800 37.780 -22.740 ;
        RECT 41.130 -22.800 41.420 -22.770 ;
        RECT 41.990 -22.800 42.310 -22.740 ;
        RECT 37.460 -22.940 42.310 -22.800 ;
        RECT 37.460 -23.000 37.780 -22.940 ;
        RECT 41.130 -23.000 41.420 -22.940 ;
        RECT 41.990 -23.000 42.310 -22.940 ;
        RECT 43.210 -22.800 43.530 -22.740 ;
        RECT 44.110 -22.800 44.400 -22.770 ;
        RECT 47.740 -22.800 48.060 -22.740 ;
        RECT 43.210 -22.940 48.060 -22.800 ;
        RECT 43.210 -23.000 43.530 -22.940 ;
        RECT 44.110 -23.000 44.400 -22.940 ;
        RECT 47.740 -23.000 48.060 -22.940 ;
        RECT 48.960 -22.800 49.280 -22.740 ;
        RECT 52.630 -22.800 52.920 -22.770 ;
        RECT 53.490 -22.800 53.810 -22.740 ;
        RECT 48.960 -22.940 53.810 -22.800 ;
        RECT 48.960 -23.000 49.280 -22.940 ;
        RECT 52.630 -23.000 52.920 -22.940 ;
        RECT 53.490 -23.000 53.810 -22.940 ;
        RECT 54.710 -22.800 55.030 -22.740 ;
        RECT 55.610 -22.800 55.900 -22.770 ;
        RECT 59.240 -22.800 59.560 -22.740 ;
        RECT 54.710 -22.940 59.560 -22.800 ;
        RECT 54.710 -23.000 55.030 -22.940 ;
        RECT 55.610 -23.000 55.900 -22.940 ;
        RECT 59.240 -23.000 59.560 -22.940 ;
        RECT 60.460 -22.800 60.780 -22.740 ;
        RECT 64.130 -22.800 64.420 -22.770 ;
        RECT 64.990 -22.800 65.310 -22.740 ;
        RECT 60.460 -22.940 65.310 -22.800 ;
        RECT 60.460 -23.000 60.780 -22.940 ;
        RECT 64.130 -23.000 64.420 -22.940 ;
        RECT 64.990 -23.000 65.310 -22.940 ;
        RECT 66.210 -22.800 66.530 -22.740 ;
        RECT 67.110 -22.800 67.400 -22.770 ;
        RECT 70.740 -22.800 71.060 -22.740 ;
        RECT 66.210 -22.940 71.060 -22.800 ;
        RECT 66.210 -23.000 66.530 -22.940 ;
        RECT 67.110 -23.000 67.400 -22.940 ;
        RECT 70.740 -23.000 71.060 -22.940 ;
        RECT 71.960 -22.800 72.280 -22.740 ;
        RECT 75.630 -22.800 75.920 -22.770 ;
        RECT 76.490 -22.800 76.810 -22.740 ;
        RECT 71.960 -22.940 76.810 -22.800 ;
        RECT 71.960 -23.000 72.280 -22.940 ;
        RECT 75.630 -23.000 75.920 -22.940 ;
        RECT 76.490 -23.000 76.810 -22.940 ;
        RECT 77.710 -22.800 78.030 -22.740 ;
        RECT 78.610 -22.800 78.900 -22.770 ;
        RECT 82.240 -22.800 82.560 -22.740 ;
        RECT 77.710 -22.940 82.560 -22.800 ;
        RECT 77.710 -23.000 78.030 -22.940 ;
        RECT 78.610 -23.000 78.900 -22.940 ;
        RECT 82.240 -23.000 82.560 -22.940 ;
        RECT 83.460 -22.800 83.780 -22.740 ;
        RECT 87.130 -22.800 87.420 -22.770 ;
        RECT 87.990 -22.800 88.310 -22.740 ;
        RECT 83.460 -22.940 88.310 -22.800 ;
        RECT 83.460 -23.000 83.780 -22.940 ;
        RECT 87.130 -23.000 87.420 -22.940 ;
        RECT 87.990 -23.000 88.310 -22.940 ;
        RECT 89.210 -22.800 89.530 -22.740 ;
        RECT 90.110 -22.800 90.400 -22.770 ;
        RECT 93.740 -22.800 94.060 -22.740 ;
        RECT 89.210 -22.940 94.060 -22.800 ;
        RECT 89.210 -23.000 89.530 -22.940 ;
        RECT 90.110 -23.000 90.400 -22.940 ;
        RECT 93.740 -23.000 94.060 -22.940 ;
        RECT 5.230 -23.670 5.550 -23.410 ;
        RECT 8.060 -23.550 8.460 -23.150 ;
        RECT 10.980 -23.680 11.300 -23.420 ;
        RECT 16.730 -23.730 17.050 -23.470 ;
        RECT 19.550 -23.560 19.950 -23.160 ;
        RECT 22.480 -23.730 22.800 -23.470 ;
        RECT 28.230 -23.730 28.550 -23.470 ;
        RECT 30.980 -23.570 31.380 -23.170 ;
        RECT 33.980 -23.730 34.300 -23.470 ;
        RECT 39.730 -23.730 40.050 -23.470 ;
        RECT 42.550 -23.580 42.950 -23.180 ;
        RECT 45.480 -23.730 45.800 -23.470 ;
        RECT 51.230 -23.730 51.550 -23.470 ;
        RECT 53.950 -23.560 54.350 -23.160 ;
        RECT 56.980 -23.730 57.300 -23.470 ;
        RECT 62.730 -23.730 63.050 -23.470 ;
        RECT 65.630 -23.560 66.030 -23.160 ;
        RECT 68.480 -23.730 68.800 -23.470 ;
        RECT 74.230 -23.730 74.550 -23.470 ;
        RECT 77.080 -23.560 77.480 -23.160 ;
        RECT 79.980 -23.730 80.300 -23.470 ;
        RECT 85.730 -23.730 86.050 -23.470 ;
        RECT 88.650 -23.540 89.050 -23.140 ;
        RECT 91.480 -23.730 91.800 -23.470 ;
        RECT 7.300 -24.540 7.700 -24.140 ;
        RECT 8.850 -24.540 9.250 -24.140 ;
        RECT 18.800 -24.540 19.200 -24.140 ;
        RECT 20.350 -24.540 20.750 -24.140 ;
        RECT 30.300 -24.540 30.700 -24.140 ;
        RECT 31.840 -24.540 32.240 -24.140 ;
        RECT 41.770 -24.540 42.170 -24.140 ;
        RECT -39.270 -24.610 -38.950 -24.580 ;
        RECT 6.620 -24.610 6.940 -24.540 ;
        RECT 43.360 -24.550 43.760 -24.150 ;
        RECT 53.290 -24.540 53.690 -24.140 ;
        RECT 54.840 -24.540 55.240 -24.140 ;
        RECT 64.800 -24.550 65.200 -24.150 ;
        RECT 66.330 -24.550 66.730 -24.150 ;
        RECT 76.310 -24.540 76.710 -24.140 ;
        RECT 77.840 -24.540 78.240 -24.140 ;
        RECT 87.800 -24.540 88.200 -24.140 ;
        RECT 89.320 -24.540 89.720 -24.130 ;
        RECT -39.270 -24.750 6.940 -24.610 ;
        RECT -39.270 -24.840 -38.950 -24.750 ;
        RECT 6.620 -24.850 6.940 -24.750 ;
        RECT 4.610 -25.310 5.010 -24.910 ;
        RECT 11.540 -25.240 11.940 -24.840 ;
        RECT 16.100 -25.230 16.500 -24.830 ;
        RECT 23.030 -25.280 23.430 -24.880 ;
        RECT 27.620 -25.290 28.020 -24.890 ;
        RECT 34.540 -25.270 34.940 -24.870 ;
        RECT 39.120 -25.290 39.520 -24.890 ;
        RECT 46.030 -25.310 46.430 -24.910 ;
        RECT 50.610 -25.250 51.010 -24.850 ;
        RECT 57.540 -25.270 57.940 -24.870 ;
        RECT 62.110 -25.230 62.510 -24.830 ;
        RECT 69.030 -25.270 69.430 -24.870 ;
        RECT 73.610 -25.270 74.010 -24.870 ;
        RECT 80.530 -25.300 80.930 -24.900 ;
        RECT 85.110 -25.290 85.510 -24.890 ;
        RECT 92.030 -25.250 92.390 -24.870 ;
        RECT -27.470 -25.450 -27.150 -25.400 ;
        RECT 9.630 -25.450 9.910 -25.400 ;
        RECT -27.470 -25.620 9.910 -25.450 ;
        RECT -27.470 -25.660 -27.150 -25.620 ;
        RECT 9.630 -25.690 9.910 -25.620 ;
        RECT 90.120 -25.420 90.410 -25.400 ;
        RECT 135.290 -25.420 135.610 -25.370 ;
        RECT 90.120 -25.590 135.610 -25.420 ;
        RECT 90.120 -25.630 90.410 -25.590 ;
        RECT 135.290 -25.630 135.610 -25.590 ;
        RECT 87.120 -25.920 87.410 -25.900 ;
        RECT 125.860 -25.920 126.120 -25.840 ;
        RECT -15.680 -26.080 -15.360 -26.030 ;
        RECT 18.120 -26.080 18.410 -26.020 ;
        RECT -15.680 -26.250 18.410 -26.080 ;
        RECT 87.120 -26.090 126.120 -25.920 ;
        RECT 87.120 -26.130 87.410 -26.090 ;
        RECT 125.860 -26.160 126.120 -26.090 ;
        RECT -15.680 -26.290 -15.360 -26.250 ;
        RECT 18.120 -26.310 18.410 -26.250 ;
        RECT 78.620 -26.420 78.910 -26.400 ;
        RECT 114.230 -26.420 114.490 -26.340 ;
        RECT 78.620 -26.590 114.490 -26.420 ;
        RECT 78.620 -26.630 78.910 -26.590 ;
        RECT 114.230 -26.660 114.490 -26.590 ;
        RECT -3.900 -26.830 -3.580 -26.780 ;
        RECT 21.120 -26.830 21.410 -26.810 ;
        RECT -3.900 -27.000 21.410 -26.830 ;
        RECT -3.900 -27.040 -3.580 -27.000 ;
        RECT 21.120 -27.040 21.410 -27.000 ;
        RECT 75.620 -27.050 75.910 -27.030 ;
        RECT 102.100 -27.050 102.360 -26.970 ;
        RECT 75.620 -27.220 102.360 -27.050 ;
        RECT 75.620 -27.260 75.910 -27.220 ;
        RECT 102.100 -27.290 102.360 -27.220 ;
        RECT 8.080 -27.540 8.400 -27.490 ;
        RECT 29.620 -27.540 29.910 -27.520 ;
        RECT 8.080 -27.710 29.910 -27.540 ;
        RECT 8.080 -27.750 8.400 -27.710 ;
        RECT 29.620 -27.750 29.910 -27.710 ;
        RECT 67.150 -27.680 67.380 -27.630 ;
        RECT 90.360 -27.680 90.620 -27.600 ;
        RECT 67.150 -27.850 90.620 -27.680 ;
        RECT 67.150 -27.920 67.380 -27.850 ;
        RECT 90.360 -27.920 90.620 -27.850 ;
        RECT 19.750 -28.340 20.070 -28.290 ;
        RECT 32.620 -28.340 32.910 -28.320 ;
        RECT 19.750 -28.510 32.910 -28.340 ;
        RECT 19.750 -28.550 20.070 -28.510 ;
        RECT 32.620 -28.550 32.910 -28.510 ;
        RECT 64.120 -28.400 64.410 -28.380 ;
        RECT 78.450 -28.400 78.770 -28.350 ;
        RECT 64.120 -28.570 78.770 -28.400 ;
        RECT 64.120 -28.610 64.410 -28.570 ;
        RECT 78.450 -28.610 78.770 -28.570 ;
        RECT 31.370 -29.180 31.630 -29.100 ;
        RECT 41.120 -29.180 41.410 -29.160 ;
        RECT 31.370 -29.350 41.410 -29.180 ;
        RECT 31.370 -29.420 31.630 -29.350 ;
        RECT 41.120 -29.390 41.410 -29.350 ;
        RECT 55.620 -29.200 55.910 -29.180 ;
        RECT 66.430 -29.200 66.750 -29.150 ;
        RECT 55.620 -29.370 66.750 -29.200 ;
        RECT 55.620 -29.410 55.910 -29.370 ;
        RECT 66.430 -29.410 66.750 -29.370 ;
        RECT 43.080 -29.890 43.400 -29.840 ;
        RECT 44.120 -29.890 44.410 -29.870 ;
        RECT 43.080 -30.060 44.410 -29.890 ;
        RECT 43.080 -30.100 43.400 -30.060 ;
        RECT 44.120 -30.100 44.410 -30.060 ;
        RECT 52.620 -30.070 52.910 -30.050 ;
        RECT 54.930 -30.070 55.250 -30.020 ;
        RECT 52.620 -30.240 55.250 -30.070 ;
        RECT 52.620 -30.280 52.910 -30.240 ;
        RECT 54.930 -30.280 55.250 -30.240 ;
        RECT -39.910 -31.310 -39.590 -31.250 ;
        RECT -37.240 -31.290 -37.010 -31.260 ;
        RECT -33.190 -31.290 -32.960 -31.260 ;
        RECT -25.740 -31.290 -25.510 -31.260 ;
        RECT -21.690 -31.290 -21.460 -31.260 ;
        RECT -13.920 -31.290 -13.690 -31.260 ;
        RECT -9.870 -31.290 -9.640 -31.260 ;
        RECT -2.110 -31.290 -1.880 -31.260 ;
        RECT 1.940 -31.290 2.170 -31.260 ;
        RECT 9.700 -31.290 9.930 -31.260 ;
        RECT 13.750 -31.290 13.980 -31.260 ;
        RECT 21.520 -31.290 21.750 -31.260 ;
        RECT 25.570 -31.290 25.800 -31.260 ;
        RECT 33.340 -31.290 33.570 -31.260 ;
        RECT 37.390 -31.290 37.620 -31.260 ;
        RECT 45.160 -31.290 45.390 -31.260 ;
        RECT 49.210 -31.290 49.440 -31.260 ;
        RECT 56.980 -31.290 57.210 -31.260 ;
        RECT 61.030 -31.290 61.260 -31.260 ;
        RECT 68.800 -31.290 69.030 -31.260 ;
        RECT 72.850 -31.290 73.080 -31.260 ;
        RECT 80.620 -31.290 80.850 -31.260 ;
        RECT 84.670 -31.290 84.900 -31.260 ;
        RECT 92.460 -31.290 92.690 -31.260 ;
        RECT 96.510 -31.290 96.740 -31.260 ;
        RECT 104.300 -31.290 104.530 -31.260 ;
        RECT 108.350 -31.290 108.580 -31.260 ;
        RECT 116.170 -31.290 116.400 -31.260 ;
        RECT 120.220 -31.290 120.450 -31.260 ;
        RECT 128.040 -31.290 128.270 -31.260 ;
        RECT 132.090 -31.290 132.320 -31.260 ;
        RECT 137.050 -31.290 137.280 -31.260 ;
        RECT 141.100 -31.290 141.330 -31.260 ;
        RECT -37.290 -31.310 -36.960 -31.290 ;
        RECT -33.240 -31.310 -32.910 -31.290 ;
        RECT -25.790 -31.310 -25.460 -31.290 ;
        RECT -21.740 -31.310 -21.410 -31.290 ;
        RECT -13.970 -31.310 -13.640 -31.290 ;
        RECT -9.920 -31.310 -9.590 -31.290 ;
        RECT -2.160 -31.310 -1.830 -31.290 ;
        RECT 1.890 -31.310 2.220 -31.290 ;
        RECT 9.650 -31.310 9.980 -31.290 ;
        RECT 13.700 -31.310 14.030 -31.290 ;
        RECT 21.470 -31.310 21.800 -31.290 ;
        RECT 25.520 -31.310 25.850 -31.290 ;
        RECT 33.290 -31.310 33.620 -31.290 ;
        RECT 37.340 -31.310 37.670 -31.290 ;
        RECT 45.110 -31.310 45.440 -31.290 ;
        RECT 49.160 -31.310 49.490 -31.290 ;
        RECT 56.930 -31.310 57.260 -31.290 ;
        RECT 60.980 -31.310 61.310 -31.290 ;
        RECT 68.750 -31.310 69.080 -31.290 ;
        RECT 72.800 -31.310 73.130 -31.290 ;
        RECT 80.570 -31.310 80.900 -31.290 ;
        RECT 84.620 -31.310 84.950 -31.290 ;
        RECT 92.410 -31.310 92.740 -31.290 ;
        RECT 96.460 -31.310 96.790 -31.290 ;
        RECT 104.250 -31.310 104.580 -31.290 ;
        RECT 108.300 -31.310 108.630 -31.290 ;
        RECT 116.120 -31.310 116.450 -31.290 ;
        RECT 120.170 -31.310 120.500 -31.290 ;
        RECT 127.990 -31.310 128.320 -31.290 ;
        RECT 132.040 -31.310 132.370 -31.290 ;
        RECT 137.000 -31.310 137.330 -31.290 ;
        RECT 141.050 -31.310 141.380 -31.290 ;
        RECT -39.910 -31.450 142.470 -31.310 ;
        RECT -39.910 -31.510 -39.590 -31.450 ;
        RECT -37.290 -31.460 -36.960 -31.450 ;
        RECT -33.240 -31.460 -32.910 -31.450 ;
        RECT -25.790 -31.460 -25.460 -31.450 ;
        RECT -21.740 -31.460 -21.410 -31.450 ;
        RECT -13.970 -31.460 -13.640 -31.450 ;
        RECT -9.920 -31.460 -9.590 -31.450 ;
        RECT -2.160 -31.460 -1.830 -31.450 ;
        RECT 1.890 -31.460 2.220 -31.450 ;
        RECT 9.650 -31.460 9.980 -31.450 ;
        RECT 13.700 -31.460 14.030 -31.450 ;
        RECT 21.470 -31.460 21.800 -31.450 ;
        RECT 25.520 -31.460 25.850 -31.450 ;
        RECT 33.290 -31.460 33.620 -31.450 ;
        RECT 37.340 -31.460 37.670 -31.450 ;
        RECT 45.110 -31.460 45.440 -31.450 ;
        RECT 49.160 -31.460 49.490 -31.450 ;
        RECT 56.930 -31.460 57.260 -31.450 ;
        RECT 60.980 -31.460 61.310 -31.450 ;
        RECT 68.750 -31.460 69.080 -31.450 ;
        RECT 72.800 -31.460 73.130 -31.450 ;
        RECT 80.570 -31.460 80.900 -31.450 ;
        RECT 84.620 -31.460 84.950 -31.450 ;
        RECT 92.410 -31.460 92.740 -31.450 ;
        RECT 96.460 -31.460 96.790 -31.450 ;
        RECT 104.250 -31.460 104.580 -31.450 ;
        RECT 108.300 -31.460 108.630 -31.450 ;
        RECT 116.120 -31.460 116.450 -31.450 ;
        RECT 120.170 -31.460 120.500 -31.450 ;
        RECT 127.990 -31.460 128.320 -31.450 ;
        RECT 132.040 -31.460 132.370 -31.450 ;
        RECT 137.000 -31.460 137.330 -31.450 ;
        RECT 141.050 -31.460 141.380 -31.450 ;
        RECT -37.240 -31.490 -37.010 -31.460 ;
        RECT -33.190 -31.490 -32.960 -31.460 ;
        RECT -25.740 -31.490 -25.510 -31.460 ;
        RECT -21.690 -31.490 -21.460 -31.460 ;
        RECT -13.920 -31.490 -13.690 -31.460 ;
        RECT -9.870 -31.490 -9.640 -31.460 ;
        RECT -2.110 -31.490 -1.880 -31.460 ;
        RECT 1.940 -31.490 2.170 -31.460 ;
        RECT 9.700 -31.490 9.930 -31.460 ;
        RECT 13.750 -31.490 13.980 -31.460 ;
        RECT 21.520 -31.490 21.750 -31.460 ;
        RECT 25.570 -31.490 25.800 -31.460 ;
        RECT 33.340 -31.490 33.570 -31.460 ;
        RECT 37.390 -31.490 37.620 -31.460 ;
        RECT 45.160 -31.490 45.390 -31.460 ;
        RECT 49.210 -31.490 49.440 -31.460 ;
        RECT 56.980 -31.490 57.210 -31.460 ;
        RECT 61.030 -31.490 61.260 -31.460 ;
        RECT 68.800 -31.490 69.030 -31.460 ;
        RECT 72.850 -31.490 73.080 -31.460 ;
        RECT 80.620 -31.490 80.850 -31.460 ;
        RECT 84.670 -31.490 84.900 -31.460 ;
        RECT 92.460 -31.490 92.690 -31.460 ;
        RECT 96.510 -31.490 96.740 -31.460 ;
        RECT 104.300 -31.490 104.530 -31.460 ;
        RECT 108.350 -31.490 108.580 -31.460 ;
        RECT 116.170 -31.490 116.400 -31.460 ;
        RECT 120.220 -31.490 120.450 -31.460 ;
        RECT 128.040 -31.490 128.270 -31.460 ;
        RECT 132.090 -31.490 132.320 -31.460 ;
        RECT 137.050 -31.490 137.280 -31.460 ;
        RECT 141.100 -31.490 141.330 -31.460 ;
        RECT -37.000 -33.670 -36.750 -33.560 ;
        RECT -35.250 -33.660 -34.930 -33.580 ;
        RECT -33.460 -33.660 -33.210 -33.570 ;
        RECT -32.350 -33.660 -32.060 -33.610 ;
        RECT -35.250 -33.670 -32.060 -33.660 ;
        RECT -37.000 -33.800 -32.060 -33.670 ;
        RECT -37.000 -33.810 -34.930 -33.800 ;
        RECT -37.000 -33.920 -36.750 -33.810 ;
        RECT -35.250 -33.900 -34.930 -33.810 ;
        RECT -33.460 -33.890 -33.210 -33.800 ;
        RECT -32.350 -33.840 -32.060 -33.800 ;
        RECT -25.500 -33.670 -25.250 -33.560 ;
        RECT -23.750 -33.660 -23.430 -33.580 ;
        RECT -21.960 -33.660 -21.710 -33.570 ;
        RECT -20.850 -33.660 -20.560 -33.610 ;
        RECT -23.750 -33.670 -20.560 -33.660 ;
        RECT -25.500 -33.800 -20.560 -33.670 ;
        RECT -25.500 -33.810 -23.430 -33.800 ;
        RECT -25.500 -33.920 -25.250 -33.810 ;
        RECT -23.750 -33.900 -23.430 -33.810 ;
        RECT -21.960 -33.890 -21.710 -33.800 ;
        RECT -20.850 -33.840 -20.560 -33.800 ;
        RECT -13.680 -33.670 -13.430 -33.560 ;
        RECT -11.930 -33.660 -11.610 -33.580 ;
        RECT -10.140 -33.660 -9.890 -33.570 ;
        RECT -9.030 -33.660 -8.740 -33.610 ;
        RECT -11.930 -33.670 -8.740 -33.660 ;
        RECT -13.680 -33.800 -8.740 -33.670 ;
        RECT -13.680 -33.810 -11.610 -33.800 ;
        RECT -13.680 -33.920 -13.430 -33.810 ;
        RECT -11.930 -33.900 -11.610 -33.810 ;
        RECT -10.140 -33.890 -9.890 -33.800 ;
        RECT -9.030 -33.840 -8.740 -33.800 ;
        RECT -1.870 -33.670 -1.620 -33.560 ;
        RECT -0.120 -33.660 0.200 -33.580 ;
        RECT 1.670 -33.660 1.920 -33.570 ;
        RECT 2.780 -33.660 3.070 -33.610 ;
        RECT -0.120 -33.670 3.070 -33.660 ;
        RECT -1.870 -33.800 3.070 -33.670 ;
        RECT -1.870 -33.810 0.200 -33.800 ;
        RECT -1.870 -33.920 -1.620 -33.810 ;
        RECT -0.120 -33.900 0.200 -33.810 ;
        RECT 1.670 -33.890 1.920 -33.800 ;
        RECT 2.780 -33.840 3.070 -33.800 ;
        RECT 9.940 -33.670 10.190 -33.560 ;
        RECT 11.690 -33.660 12.010 -33.580 ;
        RECT 13.480 -33.660 13.730 -33.570 ;
        RECT 14.590 -33.660 14.880 -33.610 ;
        RECT 11.690 -33.670 14.880 -33.660 ;
        RECT 9.940 -33.800 14.880 -33.670 ;
        RECT 9.940 -33.810 12.010 -33.800 ;
        RECT 9.940 -33.920 10.190 -33.810 ;
        RECT 11.690 -33.900 12.010 -33.810 ;
        RECT 13.480 -33.890 13.730 -33.800 ;
        RECT 14.590 -33.840 14.880 -33.800 ;
        RECT 21.760 -33.670 22.010 -33.560 ;
        RECT 23.510 -33.660 23.830 -33.580 ;
        RECT 25.300 -33.660 25.550 -33.570 ;
        RECT 26.410 -33.660 26.700 -33.610 ;
        RECT 23.510 -33.670 26.700 -33.660 ;
        RECT 21.760 -33.800 26.700 -33.670 ;
        RECT 21.760 -33.810 23.830 -33.800 ;
        RECT 21.760 -33.920 22.010 -33.810 ;
        RECT 23.510 -33.900 23.830 -33.810 ;
        RECT 25.300 -33.890 25.550 -33.800 ;
        RECT 26.410 -33.840 26.700 -33.800 ;
        RECT 33.580 -33.670 33.830 -33.560 ;
        RECT 35.330 -33.660 35.650 -33.580 ;
        RECT 37.120 -33.660 37.370 -33.570 ;
        RECT 38.230 -33.660 38.520 -33.610 ;
        RECT 35.330 -33.670 38.520 -33.660 ;
        RECT 33.580 -33.800 38.520 -33.670 ;
        RECT 33.580 -33.810 35.650 -33.800 ;
        RECT 33.580 -33.920 33.830 -33.810 ;
        RECT 35.330 -33.900 35.650 -33.810 ;
        RECT 37.120 -33.890 37.370 -33.800 ;
        RECT 38.230 -33.840 38.520 -33.800 ;
        RECT 45.400 -33.670 45.650 -33.560 ;
        RECT 47.150 -33.660 47.470 -33.580 ;
        RECT 48.940 -33.660 49.190 -33.570 ;
        RECT 50.050 -33.660 50.340 -33.610 ;
        RECT 47.150 -33.670 50.340 -33.660 ;
        RECT 45.400 -33.800 50.340 -33.670 ;
        RECT 45.400 -33.810 47.470 -33.800 ;
        RECT 45.400 -33.920 45.650 -33.810 ;
        RECT 47.150 -33.900 47.470 -33.810 ;
        RECT 48.940 -33.890 49.190 -33.800 ;
        RECT 50.050 -33.840 50.340 -33.800 ;
        RECT 57.220 -33.670 57.470 -33.560 ;
        RECT 58.970 -33.660 59.290 -33.580 ;
        RECT 60.760 -33.660 61.010 -33.570 ;
        RECT 61.870 -33.660 62.160 -33.610 ;
        RECT 58.970 -33.670 62.160 -33.660 ;
        RECT 57.220 -33.800 62.160 -33.670 ;
        RECT 57.220 -33.810 59.290 -33.800 ;
        RECT 57.220 -33.920 57.470 -33.810 ;
        RECT 58.970 -33.900 59.290 -33.810 ;
        RECT 60.760 -33.890 61.010 -33.800 ;
        RECT 61.870 -33.840 62.160 -33.800 ;
        RECT 69.040 -33.670 69.290 -33.560 ;
        RECT 70.790 -33.660 71.110 -33.580 ;
        RECT 72.580 -33.660 72.830 -33.570 ;
        RECT 73.690 -33.660 73.980 -33.610 ;
        RECT 70.790 -33.670 73.980 -33.660 ;
        RECT 69.040 -33.800 73.980 -33.670 ;
        RECT 69.040 -33.810 71.110 -33.800 ;
        RECT 69.040 -33.920 69.290 -33.810 ;
        RECT 70.790 -33.900 71.110 -33.810 ;
        RECT 72.580 -33.890 72.830 -33.800 ;
        RECT 73.690 -33.840 73.980 -33.800 ;
        RECT 80.860 -33.670 81.110 -33.560 ;
        RECT 82.610 -33.660 82.930 -33.580 ;
        RECT 84.400 -33.660 84.650 -33.570 ;
        RECT 85.510 -33.660 85.800 -33.610 ;
        RECT 82.610 -33.670 85.800 -33.660 ;
        RECT 80.860 -33.800 85.800 -33.670 ;
        RECT 80.860 -33.810 82.930 -33.800 ;
        RECT 80.860 -33.920 81.110 -33.810 ;
        RECT 82.610 -33.900 82.930 -33.810 ;
        RECT 84.400 -33.890 84.650 -33.800 ;
        RECT 85.510 -33.840 85.800 -33.800 ;
        RECT 92.700 -33.670 92.950 -33.560 ;
        RECT 94.450 -33.660 94.770 -33.580 ;
        RECT 96.240 -33.660 96.490 -33.570 ;
        RECT 97.350 -33.660 97.640 -33.610 ;
        RECT 94.450 -33.670 97.640 -33.660 ;
        RECT 92.700 -33.800 97.640 -33.670 ;
        RECT 92.700 -33.810 94.770 -33.800 ;
        RECT 92.700 -33.920 92.950 -33.810 ;
        RECT 94.450 -33.900 94.770 -33.810 ;
        RECT 96.240 -33.890 96.490 -33.800 ;
        RECT 97.350 -33.840 97.640 -33.800 ;
        RECT 104.540 -33.670 104.790 -33.560 ;
        RECT 106.290 -33.660 106.610 -33.580 ;
        RECT 108.080 -33.660 108.330 -33.570 ;
        RECT 109.190 -33.660 109.480 -33.610 ;
        RECT 106.290 -33.670 109.480 -33.660 ;
        RECT 104.540 -33.800 109.480 -33.670 ;
        RECT 104.540 -33.810 106.610 -33.800 ;
        RECT 104.540 -33.920 104.790 -33.810 ;
        RECT 106.290 -33.900 106.610 -33.810 ;
        RECT 108.080 -33.890 108.330 -33.800 ;
        RECT 109.190 -33.840 109.480 -33.800 ;
        RECT 116.410 -33.670 116.660 -33.560 ;
        RECT 118.160 -33.660 118.480 -33.580 ;
        RECT 119.950 -33.660 120.200 -33.570 ;
        RECT 121.060 -33.660 121.350 -33.610 ;
        RECT 118.160 -33.670 121.350 -33.660 ;
        RECT 116.410 -33.800 121.350 -33.670 ;
        RECT 116.410 -33.810 118.480 -33.800 ;
        RECT 116.410 -33.920 116.660 -33.810 ;
        RECT 118.160 -33.900 118.480 -33.810 ;
        RECT 119.950 -33.890 120.200 -33.800 ;
        RECT 121.060 -33.840 121.350 -33.800 ;
        RECT 128.280 -33.670 128.530 -33.560 ;
        RECT 130.030 -33.660 130.350 -33.580 ;
        RECT 131.820 -33.660 132.070 -33.570 ;
        RECT 132.930 -33.660 133.220 -33.610 ;
        RECT 130.030 -33.670 133.220 -33.660 ;
        RECT 128.280 -33.800 133.220 -33.670 ;
        RECT 128.280 -33.810 130.350 -33.800 ;
        RECT 128.280 -33.920 128.530 -33.810 ;
        RECT 130.030 -33.900 130.350 -33.810 ;
        RECT 131.820 -33.890 132.070 -33.800 ;
        RECT 132.930 -33.840 133.220 -33.800 ;
        RECT 137.290 -33.670 137.540 -33.560 ;
        RECT 139.040 -33.660 139.360 -33.580 ;
        RECT 140.830 -33.660 141.080 -33.570 ;
        RECT 141.940 -33.660 142.230 -33.610 ;
        RECT 139.040 -33.670 142.230 -33.660 ;
        RECT 137.290 -33.800 142.230 -33.670 ;
        RECT 137.290 -33.810 139.360 -33.800 ;
        RECT 137.290 -33.920 137.540 -33.810 ;
        RECT 139.040 -33.900 139.360 -33.810 ;
        RECT 140.830 -33.890 141.080 -33.800 ;
        RECT 141.940 -33.840 142.230 -33.800 ;
        RECT -36.600 -35.900 -36.310 -35.830 ;
        RECT -31.510 -35.900 -31.190 -35.840 ;
        RECT -36.600 -36.040 -31.190 -35.900 ;
        RECT -36.600 -36.120 -36.310 -36.040 ;
        RECT -31.510 -36.100 -31.190 -36.040 ;
        RECT -24.870 -35.900 -24.580 -35.830 ;
        RECT -19.960 -35.900 -19.640 -35.840 ;
        RECT -24.870 -36.040 -19.640 -35.900 ;
        RECT -24.870 -36.120 -24.580 -36.040 ;
        RECT -19.960 -36.100 -19.640 -36.040 ;
        RECT -13.120 -35.900 -12.890 -35.830 ;
        RECT -8.270 -35.900 -7.950 -35.840 ;
        RECT -13.120 -36.040 -7.950 -35.900 ;
        RECT -13.120 -36.120 -12.890 -36.040 ;
        RECT -8.270 -36.100 -7.950 -36.040 ;
        RECT -1.340 -35.900 -1.050 -35.830 ;
        RECT 3.640 -35.900 3.960 -35.840 ;
        RECT -1.340 -36.040 3.960 -35.900 ;
        RECT -1.340 -36.120 -1.050 -36.040 ;
        RECT 3.640 -36.100 3.960 -36.040 ;
        RECT 10.520 -35.900 10.810 -35.830 ;
        RECT 15.410 -35.900 15.730 -35.840 ;
        RECT 10.520 -36.040 15.730 -35.900 ;
        RECT 10.520 -36.120 10.810 -36.040 ;
        RECT 15.410 -36.100 15.730 -36.040 ;
        RECT 22.360 -35.900 22.650 -35.830 ;
        RECT 27.180 -35.900 27.500 -35.840 ;
        RECT 22.360 -36.040 27.500 -35.900 ;
        RECT 22.360 -36.120 22.650 -36.040 ;
        RECT 27.180 -36.100 27.500 -36.040 ;
        RECT 34.040 -35.900 34.330 -35.830 ;
        RECT 39.000 -35.900 39.320 -35.840 ;
        RECT 34.040 -36.040 39.320 -35.900 ;
        RECT 34.040 -36.120 34.330 -36.040 ;
        RECT 39.000 -36.100 39.320 -36.040 ;
        RECT 45.930 -35.900 46.220 -35.830 ;
        RECT 50.860 -35.900 51.180 -35.840 ;
        RECT 45.930 -36.040 51.180 -35.900 ;
        RECT 45.930 -36.120 46.220 -36.040 ;
        RECT 50.860 -36.100 51.180 -36.040 ;
        RECT 57.710 -35.900 58.000 -35.830 ;
        RECT 62.650 -35.900 62.970 -35.840 ;
        RECT 57.710 -36.040 62.970 -35.900 ;
        RECT 57.710 -36.120 58.000 -36.040 ;
        RECT 62.650 -36.100 62.970 -36.040 ;
        RECT 69.600 -35.900 69.890 -35.830 ;
        RECT 74.530 -35.900 74.850 -35.840 ;
        RECT 69.600 -36.040 74.850 -35.900 ;
        RECT 69.600 -36.120 69.890 -36.040 ;
        RECT 74.530 -36.100 74.850 -36.040 ;
        RECT 81.260 -35.900 81.550 -35.830 ;
        RECT 86.260 -35.900 86.580 -35.840 ;
        RECT 81.260 -36.040 86.580 -35.900 ;
        RECT 81.260 -36.120 81.550 -36.040 ;
        RECT 86.260 -36.100 86.580 -36.040 ;
        RECT 93.280 -35.900 93.570 -35.830 ;
        RECT 98.080 -35.900 98.400 -35.840 ;
        RECT 93.280 -36.040 98.400 -35.900 ;
        RECT 93.280 -36.120 93.570 -36.040 ;
        RECT 98.080 -36.100 98.400 -36.040 ;
        RECT 105.010 -35.900 105.300 -35.830 ;
        RECT 109.970 -35.900 110.290 -35.840 ;
        RECT 105.010 -36.040 110.290 -35.900 ;
        RECT 105.010 -36.120 105.300 -36.040 ;
        RECT 109.970 -36.100 110.290 -36.040 ;
        RECT 116.730 -35.900 117.020 -35.830 ;
        RECT 121.920 -35.900 122.240 -35.840 ;
        RECT 116.730 -36.040 122.240 -35.900 ;
        RECT 116.730 -36.120 117.020 -36.040 ;
        RECT 121.920 -36.100 122.240 -36.040 ;
        RECT 128.890 -35.900 129.180 -35.830 ;
        RECT 133.680 -35.900 134.000 -35.840 ;
        RECT 128.890 -36.040 134.000 -35.900 ;
        RECT 128.890 -36.120 129.180 -36.040 ;
        RECT 133.680 -36.100 134.000 -36.040 ;
        RECT 137.910 -35.900 138.200 -35.830 ;
        RECT 142.720 -35.900 143.040 -35.840 ;
        RECT 137.910 -36.040 143.040 -35.900 ;
        RECT 137.910 -36.120 138.200 -36.040 ;
        RECT 142.720 -36.100 143.040 -36.040 ;
        RECT -40.570 -36.340 -40.250 -36.280 ;
        RECT -36.790 -36.340 -36.460 -36.290 ;
        RECT -33.720 -36.340 -33.390 -36.280 ;
        RECT -25.290 -36.340 -24.960 -36.290 ;
        RECT -22.220 -36.340 -21.890 -36.280 ;
        RECT -13.470 -36.340 -13.140 -36.290 ;
        RECT -10.400 -36.340 -10.070 -36.280 ;
        RECT -1.660 -36.340 -1.330 -36.290 ;
        RECT 1.410 -36.340 1.740 -36.280 ;
        RECT 10.150 -36.340 10.480 -36.290 ;
        RECT 13.220 -36.340 13.550 -36.280 ;
        RECT 21.970 -36.340 22.300 -36.290 ;
        RECT 25.040 -36.340 25.370 -36.280 ;
        RECT 33.790 -36.340 34.120 -36.290 ;
        RECT 36.860 -36.340 37.190 -36.280 ;
        RECT 45.610 -36.340 45.940 -36.290 ;
        RECT 48.680 -36.340 49.010 -36.280 ;
        RECT 57.430 -36.340 57.760 -36.290 ;
        RECT 60.500 -36.340 60.830 -36.280 ;
        RECT 69.250 -36.340 69.580 -36.290 ;
        RECT 72.320 -36.340 72.650 -36.280 ;
        RECT 81.070 -36.340 81.400 -36.290 ;
        RECT 84.140 -36.340 84.470 -36.280 ;
        RECT 92.910 -36.340 93.240 -36.290 ;
        RECT 95.980 -36.340 96.310 -36.280 ;
        RECT 104.750 -36.340 105.080 -36.290 ;
        RECT 107.820 -36.340 108.150 -36.280 ;
        RECT 116.620 -36.340 116.950 -36.290 ;
        RECT 119.690 -36.340 120.020 -36.280 ;
        RECT 128.490 -36.340 128.820 -36.290 ;
        RECT 131.560 -36.340 131.890 -36.280 ;
        RECT 137.500 -36.340 137.830 -36.290 ;
        RECT 140.570 -36.340 140.900 -36.280 ;
        RECT -40.570 -36.480 142.470 -36.340 ;
        RECT -40.570 -36.540 -40.250 -36.480 ;
        RECT -36.790 -36.530 -36.460 -36.480 ;
        RECT -33.720 -36.520 -33.390 -36.480 ;
        RECT -25.290 -36.530 -24.960 -36.480 ;
        RECT -22.220 -36.520 -21.890 -36.480 ;
        RECT -13.470 -36.530 -13.140 -36.480 ;
        RECT -10.400 -36.520 -10.070 -36.480 ;
        RECT -1.660 -36.530 -1.330 -36.480 ;
        RECT 1.410 -36.520 1.740 -36.480 ;
        RECT 10.150 -36.530 10.480 -36.480 ;
        RECT 13.220 -36.520 13.550 -36.480 ;
        RECT 21.970 -36.530 22.300 -36.480 ;
        RECT 25.040 -36.520 25.370 -36.480 ;
        RECT 33.790 -36.530 34.120 -36.480 ;
        RECT 36.860 -36.520 37.190 -36.480 ;
        RECT 45.610 -36.530 45.940 -36.480 ;
        RECT 48.680 -36.520 49.010 -36.480 ;
        RECT 57.430 -36.530 57.760 -36.480 ;
        RECT 60.500 -36.520 60.830 -36.480 ;
        RECT 69.250 -36.530 69.580 -36.480 ;
        RECT 72.320 -36.520 72.650 -36.480 ;
        RECT 81.070 -36.530 81.400 -36.480 ;
        RECT 84.140 -36.520 84.470 -36.480 ;
        RECT 92.910 -36.530 93.240 -36.480 ;
        RECT 95.980 -36.520 96.310 -36.480 ;
        RECT 104.750 -36.530 105.080 -36.480 ;
        RECT 107.820 -36.520 108.150 -36.480 ;
        RECT 116.620 -36.530 116.950 -36.480 ;
        RECT 119.690 -36.520 120.020 -36.480 ;
        RECT 128.490 -36.530 128.820 -36.480 ;
        RECT 131.560 -36.520 131.890 -36.480 ;
        RECT 137.500 -36.530 137.830 -36.480 ;
        RECT 140.570 -36.520 140.900 -36.480 ;
        RECT -41.230 -36.740 -40.910 -36.680 ;
        RECT -37.860 -36.710 -37.570 -36.680 ;
        RECT -37.900 -36.740 -37.570 -36.710 ;
        RECT -32.640 -36.730 -32.350 -36.700 ;
        RECT -26.360 -36.710 -26.070 -36.680 ;
        RECT -32.640 -36.740 -32.310 -36.730 ;
        RECT -26.400 -36.740 -26.070 -36.710 ;
        RECT -21.140 -36.730 -20.850 -36.700 ;
        RECT -14.540 -36.710 -14.250 -36.680 ;
        RECT -21.140 -36.740 -20.810 -36.730 ;
        RECT -14.580 -36.740 -14.250 -36.710 ;
        RECT -9.320 -36.730 -9.030 -36.700 ;
        RECT -2.730 -36.710 -2.440 -36.680 ;
        RECT -9.320 -36.740 -8.990 -36.730 ;
        RECT -2.770 -36.740 -2.440 -36.710 ;
        RECT 2.490 -36.730 2.780 -36.700 ;
        RECT 9.080 -36.710 9.370 -36.680 ;
        RECT 2.490 -36.740 2.820 -36.730 ;
        RECT 9.040 -36.740 9.370 -36.710 ;
        RECT 14.300 -36.730 14.590 -36.700 ;
        RECT 20.900 -36.710 21.190 -36.680 ;
        RECT 14.300 -36.740 14.630 -36.730 ;
        RECT 20.860 -36.740 21.190 -36.710 ;
        RECT 26.120 -36.730 26.410 -36.700 ;
        RECT 32.720 -36.710 33.010 -36.680 ;
        RECT 26.120 -36.740 26.450 -36.730 ;
        RECT 32.680 -36.740 33.010 -36.710 ;
        RECT 37.940 -36.730 38.230 -36.700 ;
        RECT 44.540 -36.710 44.830 -36.680 ;
        RECT 37.940 -36.740 38.270 -36.730 ;
        RECT 44.500 -36.740 44.830 -36.710 ;
        RECT 49.760 -36.730 50.050 -36.700 ;
        RECT 56.360 -36.710 56.650 -36.680 ;
        RECT 49.760 -36.740 50.090 -36.730 ;
        RECT 56.320 -36.740 56.650 -36.710 ;
        RECT 61.580 -36.730 61.870 -36.700 ;
        RECT 68.180 -36.710 68.470 -36.680 ;
        RECT 61.580 -36.740 61.910 -36.730 ;
        RECT 68.140 -36.740 68.470 -36.710 ;
        RECT 73.400 -36.730 73.690 -36.700 ;
        RECT 80.000 -36.710 80.290 -36.680 ;
        RECT 73.400 -36.740 73.730 -36.730 ;
        RECT 79.960 -36.740 80.290 -36.710 ;
        RECT 85.220 -36.730 85.510 -36.700 ;
        RECT 91.840 -36.710 92.130 -36.680 ;
        RECT 85.220 -36.740 85.550 -36.730 ;
        RECT 91.800 -36.740 92.130 -36.710 ;
        RECT 97.060 -36.730 97.350 -36.700 ;
        RECT 103.680 -36.710 103.970 -36.680 ;
        RECT 97.060 -36.740 97.390 -36.730 ;
        RECT 103.640 -36.740 103.970 -36.710 ;
        RECT 108.900 -36.730 109.190 -36.700 ;
        RECT 115.550 -36.710 115.840 -36.680 ;
        RECT 108.900 -36.740 109.230 -36.730 ;
        RECT 115.510 -36.740 115.840 -36.710 ;
        RECT 120.770 -36.730 121.060 -36.700 ;
        RECT 127.420 -36.710 127.710 -36.680 ;
        RECT 120.770 -36.740 121.100 -36.730 ;
        RECT 127.380 -36.740 127.710 -36.710 ;
        RECT 132.640 -36.730 132.930 -36.700 ;
        RECT 136.430 -36.710 136.720 -36.680 ;
        RECT 132.640 -36.740 132.970 -36.730 ;
        RECT 136.390 -36.740 136.720 -36.710 ;
        RECT 141.650 -36.730 141.940 -36.700 ;
        RECT 141.650 -36.740 141.980 -36.730 ;
        RECT -41.230 -36.880 142.470 -36.740 ;
        RECT -41.230 -36.940 -40.910 -36.880 ;
        RECT -37.900 -36.890 -37.570 -36.880 ;
        RECT -37.860 -36.920 -37.570 -36.890 ;
        RECT -32.640 -36.910 -32.310 -36.880 ;
        RECT -26.400 -36.890 -26.070 -36.880 ;
        RECT -32.640 -36.940 -32.350 -36.910 ;
        RECT -26.360 -36.920 -26.070 -36.890 ;
        RECT -21.140 -36.910 -20.810 -36.880 ;
        RECT -14.580 -36.890 -14.250 -36.880 ;
        RECT -21.140 -36.940 -20.850 -36.910 ;
        RECT -14.540 -36.920 -14.250 -36.890 ;
        RECT -9.320 -36.910 -8.990 -36.880 ;
        RECT -2.770 -36.890 -2.440 -36.880 ;
        RECT -9.320 -36.940 -9.030 -36.910 ;
        RECT -2.730 -36.920 -2.440 -36.890 ;
        RECT 2.490 -36.910 2.820 -36.880 ;
        RECT 9.040 -36.890 9.370 -36.880 ;
        RECT 2.490 -36.940 2.780 -36.910 ;
        RECT 9.080 -36.920 9.370 -36.890 ;
        RECT 14.300 -36.910 14.630 -36.880 ;
        RECT 20.860 -36.890 21.190 -36.880 ;
        RECT 14.300 -36.940 14.590 -36.910 ;
        RECT 20.900 -36.920 21.190 -36.890 ;
        RECT 26.120 -36.910 26.450 -36.880 ;
        RECT 32.680 -36.890 33.010 -36.880 ;
        RECT 26.120 -36.940 26.410 -36.910 ;
        RECT 32.720 -36.920 33.010 -36.890 ;
        RECT 37.940 -36.910 38.270 -36.880 ;
        RECT 44.500 -36.890 44.830 -36.880 ;
        RECT 37.940 -36.940 38.230 -36.910 ;
        RECT 44.540 -36.920 44.830 -36.890 ;
        RECT 49.760 -36.910 50.090 -36.880 ;
        RECT 56.320 -36.890 56.650 -36.880 ;
        RECT 49.760 -36.940 50.050 -36.910 ;
        RECT 56.360 -36.920 56.650 -36.890 ;
        RECT 61.580 -36.910 61.910 -36.880 ;
        RECT 68.140 -36.890 68.470 -36.880 ;
        RECT 61.580 -36.940 61.870 -36.910 ;
        RECT 68.180 -36.920 68.470 -36.890 ;
        RECT 73.400 -36.910 73.730 -36.880 ;
        RECT 79.960 -36.890 80.290 -36.880 ;
        RECT 73.400 -36.940 73.690 -36.910 ;
        RECT 80.000 -36.920 80.290 -36.890 ;
        RECT 85.220 -36.910 85.550 -36.880 ;
        RECT 91.800 -36.890 92.130 -36.880 ;
        RECT 85.220 -36.940 85.510 -36.910 ;
        RECT 91.840 -36.920 92.130 -36.890 ;
        RECT 97.060 -36.910 97.390 -36.880 ;
        RECT 103.640 -36.890 103.970 -36.880 ;
        RECT 97.060 -36.940 97.350 -36.910 ;
        RECT 103.680 -36.920 103.970 -36.890 ;
        RECT 108.900 -36.910 109.230 -36.880 ;
        RECT 115.510 -36.890 115.840 -36.880 ;
        RECT 108.900 -36.940 109.190 -36.910 ;
        RECT 115.550 -36.920 115.840 -36.890 ;
        RECT 120.770 -36.910 121.100 -36.880 ;
        RECT 127.380 -36.890 127.710 -36.880 ;
        RECT 120.770 -36.940 121.060 -36.910 ;
        RECT 127.420 -36.920 127.710 -36.890 ;
        RECT 132.640 -36.910 132.970 -36.880 ;
        RECT 136.390 -36.890 136.720 -36.880 ;
        RECT 132.640 -36.940 132.930 -36.910 ;
        RECT 136.430 -36.920 136.720 -36.890 ;
        RECT 141.650 -36.910 141.980 -36.880 ;
        RECT 141.650 -36.940 141.940 -36.910 ;
        RECT -37.940 -37.370 -37.650 -37.310 ;
        RECT -36.460 -37.370 -36.170 -37.280 ;
        RECT -37.940 -37.510 -36.170 -37.370 ;
        RECT -37.940 -37.560 -37.650 -37.510 ;
        RECT -36.460 -37.530 -36.170 -37.510 ;
        RECT -34.010 -37.340 -33.720 -37.270 ;
        RECT -32.560 -37.340 -32.270 -37.300 ;
        RECT -34.010 -37.480 -32.270 -37.340 ;
        RECT -34.010 -37.520 -33.720 -37.480 ;
        RECT -32.560 -37.550 -32.270 -37.480 ;
        RECT -26.440 -37.370 -26.150 -37.310 ;
        RECT -24.960 -37.370 -24.670 -37.280 ;
        RECT -26.440 -37.510 -24.670 -37.370 ;
        RECT -26.440 -37.560 -26.150 -37.510 ;
        RECT -24.960 -37.530 -24.670 -37.510 ;
        RECT -22.510 -37.340 -22.220 -37.270 ;
        RECT -21.060 -37.340 -20.770 -37.300 ;
        RECT -22.510 -37.480 -20.770 -37.340 ;
        RECT -22.510 -37.520 -22.220 -37.480 ;
        RECT -21.060 -37.550 -20.770 -37.480 ;
        RECT -14.620 -37.370 -14.330 -37.310 ;
        RECT -13.140 -37.370 -12.850 -37.280 ;
        RECT -14.620 -37.510 -12.850 -37.370 ;
        RECT -14.620 -37.560 -14.330 -37.510 ;
        RECT -13.140 -37.530 -12.850 -37.510 ;
        RECT -10.690 -37.340 -10.400 -37.270 ;
        RECT -9.240 -37.340 -8.950 -37.300 ;
        RECT -10.690 -37.480 -8.950 -37.340 ;
        RECT -10.690 -37.520 -10.400 -37.480 ;
        RECT -9.240 -37.550 -8.950 -37.480 ;
        RECT -2.810 -37.370 -2.520 -37.310 ;
        RECT -1.330 -37.370 -1.040 -37.280 ;
        RECT -2.810 -37.510 -1.040 -37.370 ;
        RECT -2.810 -37.560 -2.520 -37.510 ;
        RECT -1.330 -37.530 -1.040 -37.510 ;
        RECT 1.120 -37.340 1.410 -37.270 ;
        RECT 2.570 -37.340 2.860 -37.300 ;
        RECT 1.120 -37.480 2.860 -37.340 ;
        RECT 1.120 -37.520 1.410 -37.480 ;
        RECT 2.570 -37.550 2.860 -37.480 ;
        RECT 9.000 -37.370 9.290 -37.310 ;
        RECT 10.480 -37.370 10.770 -37.280 ;
        RECT 9.000 -37.510 10.770 -37.370 ;
        RECT 9.000 -37.560 9.290 -37.510 ;
        RECT 10.480 -37.530 10.770 -37.510 ;
        RECT 12.930 -37.340 13.220 -37.270 ;
        RECT 14.380 -37.340 14.670 -37.300 ;
        RECT 12.930 -37.480 14.670 -37.340 ;
        RECT 12.930 -37.520 13.220 -37.480 ;
        RECT 14.380 -37.550 14.670 -37.480 ;
        RECT 20.820 -37.370 21.110 -37.310 ;
        RECT 22.300 -37.370 22.590 -37.280 ;
        RECT 20.820 -37.510 22.590 -37.370 ;
        RECT 20.820 -37.560 21.110 -37.510 ;
        RECT 22.300 -37.530 22.590 -37.510 ;
        RECT 24.750 -37.340 25.040 -37.270 ;
        RECT 26.200 -37.340 26.490 -37.300 ;
        RECT 24.750 -37.480 26.490 -37.340 ;
        RECT 24.750 -37.520 25.040 -37.480 ;
        RECT 26.200 -37.550 26.490 -37.480 ;
        RECT 32.640 -37.370 32.930 -37.310 ;
        RECT 34.120 -37.370 34.410 -37.280 ;
        RECT 32.640 -37.510 34.410 -37.370 ;
        RECT 32.640 -37.560 32.930 -37.510 ;
        RECT 34.120 -37.530 34.410 -37.510 ;
        RECT 36.570 -37.340 36.860 -37.270 ;
        RECT 38.020 -37.340 38.310 -37.300 ;
        RECT 36.570 -37.480 38.310 -37.340 ;
        RECT 36.570 -37.520 36.860 -37.480 ;
        RECT 38.020 -37.550 38.310 -37.480 ;
        RECT 44.460 -37.370 44.750 -37.310 ;
        RECT 45.940 -37.370 46.230 -37.280 ;
        RECT 44.460 -37.510 46.230 -37.370 ;
        RECT 44.460 -37.560 44.750 -37.510 ;
        RECT 45.940 -37.530 46.230 -37.510 ;
        RECT 48.390 -37.340 48.680 -37.270 ;
        RECT 49.840 -37.340 50.130 -37.300 ;
        RECT 48.390 -37.480 50.130 -37.340 ;
        RECT 48.390 -37.520 48.680 -37.480 ;
        RECT 49.840 -37.550 50.130 -37.480 ;
        RECT 56.280 -37.370 56.570 -37.310 ;
        RECT 57.760 -37.370 58.050 -37.280 ;
        RECT 56.280 -37.510 58.050 -37.370 ;
        RECT 56.280 -37.560 56.570 -37.510 ;
        RECT 57.760 -37.530 58.050 -37.510 ;
        RECT 60.210 -37.340 60.500 -37.270 ;
        RECT 61.660 -37.340 61.950 -37.300 ;
        RECT 60.210 -37.480 61.950 -37.340 ;
        RECT 60.210 -37.520 60.500 -37.480 ;
        RECT 61.660 -37.550 61.950 -37.480 ;
        RECT 68.100 -37.370 68.390 -37.310 ;
        RECT 69.580 -37.370 69.870 -37.280 ;
        RECT 68.100 -37.510 69.870 -37.370 ;
        RECT 68.100 -37.560 68.390 -37.510 ;
        RECT 69.580 -37.530 69.870 -37.510 ;
        RECT 72.030 -37.340 72.320 -37.270 ;
        RECT 73.480 -37.340 73.770 -37.300 ;
        RECT 72.030 -37.480 73.770 -37.340 ;
        RECT 72.030 -37.520 72.320 -37.480 ;
        RECT 73.480 -37.550 73.770 -37.480 ;
        RECT 79.920 -37.370 80.210 -37.310 ;
        RECT 81.400 -37.370 81.690 -37.280 ;
        RECT 79.920 -37.510 81.690 -37.370 ;
        RECT 79.920 -37.560 80.210 -37.510 ;
        RECT 81.400 -37.530 81.690 -37.510 ;
        RECT 83.850 -37.340 84.140 -37.270 ;
        RECT 85.300 -37.340 85.590 -37.300 ;
        RECT 83.850 -37.480 85.590 -37.340 ;
        RECT 83.850 -37.520 84.140 -37.480 ;
        RECT 85.300 -37.550 85.590 -37.480 ;
        RECT 91.760 -37.370 92.050 -37.310 ;
        RECT 93.240 -37.370 93.530 -37.280 ;
        RECT 91.760 -37.510 93.530 -37.370 ;
        RECT 91.760 -37.560 92.050 -37.510 ;
        RECT 93.240 -37.530 93.530 -37.510 ;
        RECT 95.690 -37.340 95.980 -37.270 ;
        RECT 97.140 -37.340 97.430 -37.300 ;
        RECT 95.690 -37.480 97.430 -37.340 ;
        RECT 95.690 -37.520 95.980 -37.480 ;
        RECT 97.140 -37.550 97.430 -37.480 ;
        RECT 103.600 -37.370 103.890 -37.310 ;
        RECT 105.080 -37.370 105.370 -37.280 ;
        RECT 103.600 -37.510 105.370 -37.370 ;
        RECT 103.600 -37.560 103.890 -37.510 ;
        RECT 105.080 -37.530 105.370 -37.510 ;
        RECT 107.530 -37.340 107.820 -37.270 ;
        RECT 108.980 -37.340 109.270 -37.300 ;
        RECT 107.530 -37.480 109.270 -37.340 ;
        RECT 107.530 -37.520 107.820 -37.480 ;
        RECT 108.980 -37.550 109.270 -37.480 ;
        RECT 115.470 -37.370 115.760 -37.310 ;
        RECT 116.950 -37.370 117.240 -37.280 ;
        RECT 115.470 -37.510 117.240 -37.370 ;
        RECT 115.470 -37.560 115.760 -37.510 ;
        RECT 116.950 -37.530 117.240 -37.510 ;
        RECT 119.400 -37.340 119.690 -37.270 ;
        RECT 120.850 -37.340 121.140 -37.300 ;
        RECT 119.400 -37.480 121.140 -37.340 ;
        RECT 119.400 -37.520 119.690 -37.480 ;
        RECT 120.850 -37.550 121.140 -37.480 ;
        RECT 127.340 -37.370 127.630 -37.310 ;
        RECT 128.820 -37.370 129.110 -37.280 ;
        RECT 127.340 -37.510 129.110 -37.370 ;
        RECT 127.340 -37.560 127.630 -37.510 ;
        RECT 128.820 -37.530 129.110 -37.510 ;
        RECT 131.270 -37.340 131.560 -37.270 ;
        RECT 132.720 -37.340 133.010 -37.300 ;
        RECT 131.270 -37.480 133.010 -37.340 ;
        RECT 131.270 -37.520 131.560 -37.480 ;
        RECT 132.720 -37.550 133.010 -37.480 ;
        RECT 136.350 -37.370 136.640 -37.310 ;
        RECT 137.830 -37.370 138.120 -37.280 ;
        RECT 136.350 -37.510 138.120 -37.370 ;
        RECT 136.350 -37.560 136.640 -37.510 ;
        RECT 137.830 -37.530 138.120 -37.510 ;
        RECT 140.280 -37.340 140.570 -37.270 ;
        RECT 141.730 -37.340 142.020 -37.300 ;
        RECT 140.280 -37.480 142.020 -37.340 ;
        RECT 140.280 -37.520 140.570 -37.480 ;
        RECT 141.730 -37.550 142.020 -37.480 ;
        RECT -36.460 -38.040 -36.170 -37.990 ;
        RECT -35.500 -38.040 -35.210 -37.990 ;
        RECT -36.460 -38.180 -35.210 -38.040 ;
        RECT -36.460 -38.240 -36.170 -38.180 ;
        RECT -35.500 -38.240 -35.210 -38.180 ;
        RECT -24.960 -38.040 -24.670 -37.990 ;
        RECT -24.000 -38.040 -23.710 -37.990 ;
        RECT -24.960 -38.180 -23.710 -38.040 ;
        RECT -24.960 -38.240 -24.670 -38.180 ;
        RECT -24.000 -38.240 -23.710 -38.180 ;
        RECT -13.140 -38.040 -12.850 -37.990 ;
        RECT -12.180 -38.040 -11.890 -37.990 ;
        RECT -13.140 -38.180 -11.890 -38.040 ;
        RECT -13.140 -38.240 -12.850 -38.180 ;
        RECT -12.180 -38.240 -11.890 -38.180 ;
        RECT -1.330 -38.040 -1.040 -37.990 ;
        RECT -0.370 -38.040 -0.080 -37.990 ;
        RECT -1.330 -38.180 -0.080 -38.040 ;
        RECT -1.330 -38.240 -1.040 -38.180 ;
        RECT -0.370 -38.240 -0.080 -38.180 ;
        RECT 10.480 -38.040 10.770 -37.990 ;
        RECT 11.440 -38.040 11.730 -37.990 ;
        RECT 10.480 -38.180 11.730 -38.040 ;
        RECT 10.480 -38.240 10.770 -38.180 ;
        RECT 11.440 -38.240 11.730 -38.180 ;
        RECT 22.300 -38.040 22.590 -37.990 ;
        RECT 23.260 -38.040 23.550 -37.990 ;
        RECT 22.300 -38.180 23.550 -38.040 ;
        RECT 22.300 -38.240 22.590 -38.180 ;
        RECT 23.260 -38.240 23.550 -38.180 ;
        RECT 34.120 -38.040 34.410 -37.990 ;
        RECT 35.080 -38.040 35.370 -37.990 ;
        RECT 34.120 -38.180 35.370 -38.040 ;
        RECT 34.120 -38.240 34.410 -38.180 ;
        RECT 35.080 -38.240 35.370 -38.180 ;
        RECT 45.940 -38.040 46.230 -37.990 ;
        RECT 46.900 -38.040 47.190 -37.990 ;
        RECT 45.940 -38.180 47.190 -38.040 ;
        RECT 45.940 -38.240 46.230 -38.180 ;
        RECT 46.900 -38.240 47.190 -38.180 ;
        RECT 57.760 -38.040 58.050 -37.990 ;
        RECT 58.720 -38.040 59.010 -37.990 ;
        RECT 57.760 -38.180 59.010 -38.040 ;
        RECT 57.760 -38.240 58.050 -38.180 ;
        RECT 58.720 -38.240 59.010 -38.180 ;
        RECT 69.580 -38.040 69.870 -37.990 ;
        RECT 70.540 -38.040 70.830 -37.990 ;
        RECT 69.580 -38.180 70.830 -38.040 ;
        RECT 69.580 -38.240 69.870 -38.180 ;
        RECT 70.540 -38.240 70.830 -38.180 ;
        RECT 81.400 -38.040 81.690 -37.990 ;
        RECT 82.360 -38.040 82.650 -37.990 ;
        RECT 81.400 -38.180 82.650 -38.040 ;
        RECT 81.400 -38.240 81.690 -38.180 ;
        RECT 82.360 -38.240 82.650 -38.180 ;
        RECT 93.240 -38.040 93.530 -37.990 ;
        RECT 94.200 -38.040 94.490 -37.990 ;
        RECT 93.240 -38.180 94.490 -38.040 ;
        RECT 93.240 -38.240 93.530 -38.180 ;
        RECT 94.200 -38.240 94.490 -38.180 ;
        RECT 105.080 -38.040 105.370 -37.990 ;
        RECT 106.040 -38.040 106.330 -37.990 ;
        RECT 105.080 -38.180 106.330 -38.040 ;
        RECT 105.080 -38.240 105.370 -38.180 ;
        RECT 106.040 -38.240 106.330 -38.180 ;
        RECT 116.950 -38.040 117.240 -37.990 ;
        RECT 117.910 -38.040 118.200 -37.990 ;
        RECT 116.950 -38.180 118.200 -38.040 ;
        RECT 116.950 -38.240 117.240 -38.180 ;
        RECT 117.910 -38.240 118.200 -38.180 ;
        RECT 128.820 -38.040 129.110 -37.990 ;
        RECT 129.780 -38.040 130.070 -37.990 ;
        RECT 128.820 -38.180 130.070 -38.040 ;
        RECT 128.820 -38.240 129.110 -38.180 ;
        RECT 129.780 -38.240 130.070 -38.180 ;
        RECT 137.830 -38.040 138.120 -37.990 ;
        RECT 138.790 -38.040 139.080 -37.990 ;
        RECT 137.830 -38.180 139.080 -38.040 ;
        RECT 137.830 -38.240 138.120 -38.180 ;
        RECT 138.790 -38.240 139.080 -38.180 ;
        RECT -34.970 -38.850 -34.680 -38.800 ;
        RECT -34.010 -38.850 -33.720 -38.810 ;
        RECT -34.970 -38.990 -33.720 -38.850 ;
        RECT -34.970 -39.050 -34.680 -38.990 ;
        RECT -34.010 -39.060 -33.720 -38.990 ;
        RECT -23.470 -38.850 -23.180 -38.800 ;
        RECT -22.510 -38.850 -22.220 -38.810 ;
        RECT -23.470 -38.990 -22.220 -38.850 ;
        RECT -23.470 -39.050 -23.180 -38.990 ;
        RECT -22.510 -39.060 -22.220 -38.990 ;
        RECT -11.650 -38.850 -11.360 -38.800 ;
        RECT -10.690 -38.850 -10.400 -38.810 ;
        RECT -11.650 -38.990 -10.400 -38.850 ;
        RECT -11.650 -39.050 -11.360 -38.990 ;
        RECT -10.690 -39.060 -10.400 -38.990 ;
        RECT 0.160 -38.850 0.450 -38.800 ;
        RECT 1.120 -38.850 1.410 -38.810 ;
        RECT 0.160 -38.990 1.410 -38.850 ;
        RECT 0.160 -39.050 0.450 -38.990 ;
        RECT 1.120 -39.060 1.410 -38.990 ;
        RECT 11.970 -38.850 12.260 -38.800 ;
        RECT 12.930 -38.850 13.220 -38.810 ;
        RECT 11.970 -38.990 13.220 -38.850 ;
        RECT 11.970 -39.050 12.260 -38.990 ;
        RECT 12.930 -39.060 13.220 -38.990 ;
        RECT 23.790 -38.850 24.080 -38.800 ;
        RECT 24.750 -38.850 25.040 -38.810 ;
        RECT 23.790 -38.990 25.040 -38.850 ;
        RECT 23.790 -39.050 24.080 -38.990 ;
        RECT 24.750 -39.060 25.040 -38.990 ;
        RECT 35.610 -38.850 35.900 -38.800 ;
        RECT 36.570 -38.850 36.860 -38.810 ;
        RECT 35.610 -38.990 36.860 -38.850 ;
        RECT 35.610 -39.050 35.900 -38.990 ;
        RECT 36.570 -39.060 36.860 -38.990 ;
        RECT 47.430 -38.850 47.720 -38.800 ;
        RECT 48.390 -38.850 48.680 -38.810 ;
        RECT 47.430 -38.990 48.680 -38.850 ;
        RECT 47.430 -39.050 47.720 -38.990 ;
        RECT 48.390 -39.060 48.680 -38.990 ;
        RECT 59.250 -38.850 59.540 -38.800 ;
        RECT 60.210 -38.850 60.500 -38.810 ;
        RECT 59.250 -38.990 60.500 -38.850 ;
        RECT 59.250 -39.050 59.540 -38.990 ;
        RECT 60.210 -39.060 60.500 -38.990 ;
        RECT 71.070 -38.850 71.360 -38.800 ;
        RECT 72.030 -38.850 72.320 -38.810 ;
        RECT 71.070 -38.990 72.320 -38.850 ;
        RECT 71.070 -39.050 71.360 -38.990 ;
        RECT 72.030 -39.060 72.320 -38.990 ;
        RECT 82.890 -38.850 83.180 -38.800 ;
        RECT 83.850 -38.850 84.140 -38.810 ;
        RECT 82.890 -38.990 84.140 -38.850 ;
        RECT 82.890 -39.050 83.180 -38.990 ;
        RECT 83.850 -39.060 84.140 -38.990 ;
        RECT 94.730 -38.850 95.020 -38.800 ;
        RECT 95.690 -38.850 95.980 -38.810 ;
        RECT 94.730 -38.990 95.980 -38.850 ;
        RECT 94.730 -39.050 95.020 -38.990 ;
        RECT 95.690 -39.060 95.980 -38.990 ;
        RECT 106.570 -38.850 106.860 -38.800 ;
        RECT 107.530 -38.850 107.820 -38.810 ;
        RECT 106.570 -38.990 107.820 -38.850 ;
        RECT 106.570 -39.050 106.860 -38.990 ;
        RECT 107.530 -39.060 107.820 -38.990 ;
        RECT 118.440 -38.850 118.730 -38.800 ;
        RECT 119.400 -38.850 119.690 -38.810 ;
        RECT 118.440 -38.990 119.690 -38.850 ;
        RECT 118.440 -39.050 118.730 -38.990 ;
        RECT 119.400 -39.060 119.690 -38.990 ;
        RECT 130.310 -38.850 130.600 -38.800 ;
        RECT 131.270 -38.850 131.560 -38.810 ;
        RECT 130.310 -38.990 131.560 -38.850 ;
        RECT 130.310 -39.050 130.600 -38.990 ;
        RECT 131.270 -39.060 131.560 -38.990 ;
        RECT 139.320 -38.850 139.610 -38.800 ;
        RECT 140.280 -38.850 140.570 -38.810 ;
        RECT 139.320 -38.990 140.570 -38.850 ;
        RECT 139.320 -39.050 139.610 -38.990 ;
        RECT 140.280 -39.060 140.570 -38.990 ;
        RECT -38.290 -39.590 -38.000 -39.540 ;
        RECT -36.900 -39.590 -36.610 -39.540 ;
        RECT -38.290 -39.730 -36.610 -39.590 ;
        RECT -38.290 -39.790 -38.000 -39.730 ;
        RECT -36.900 -39.790 -36.610 -39.730 ;
        RECT -33.570 -39.590 -33.280 -39.530 ;
        RECT -32.210 -39.590 -31.920 -39.540 ;
        RECT -33.570 -39.730 -31.920 -39.590 ;
        RECT -33.570 -39.780 -33.280 -39.730 ;
        RECT -32.210 -39.790 -31.920 -39.730 ;
        RECT -26.790 -39.590 -26.500 -39.540 ;
        RECT -25.400 -39.590 -25.110 -39.540 ;
        RECT -26.790 -39.730 -25.110 -39.590 ;
        RECT -26.790 -39.790 -26.500 -39.730 ;
        RECT -25.400 -39.790 -25.110 -39.730 ;
        RECT -22.070 -39.590 -21.780 -39.530 ;
        RECT -20.710 -39.590 -20.420 -39.540 ;
        RECT -22.070 -39.730 -20.420 -39.590 ;
        RECT -22.070 -39.780 -21.780 -39.730 ;
        RECT -20.710 -39.790 -20.420 -39.730 ;
        RECT -14.970 -39.590 -14.680 -39.540 ;
        RECT -13.580 -39.590 -13.290 -39.540 ;
        RECT -14.970 -39.730 -13.290 -39.590 ;
        RECT -14.970 -39.790 -14.680 -39.730 ;
        RECT -13.580 -39.790 -13.290 -39.730 ;
        RECT -10.250 -39.590 -9.960 -39.530 ;
        RECT -8.890 -39.590 -8.600 -39.540 ;
        RECT -10.250 -39.730 -8.600 -39.590 ;
        RECT -10.250 -39.780 -9.960 -39.730 ;
        RECT -8.890 -39.790 -8.600 -39.730 ;
        RECT -3.160 -39.590 -2.870 -39.540 ;
        RECT -1.770 -39.590 -1.480 -39.540 ;
        RECT -3.160 -39.730 -1.480 -39.590 ;
        RECT -3.160 -39.790 -2.870 -39.730 ;
        RECT -1.770 -39.790 -1.480 -39.730 ;
        RECT 1.560 -39.590 1.850 -39.530 ;
        RECT 2.920 -39.590 3.210 -39.540 ;
        RECT 1.560 -39.730 3.210 -39.590 ;
        RECT 1.560 -39.780 1.850 -39.730 ;
        RECT 2.920 -39.790 3.210 -39.730 ;
        RECT 8.650 -39.590 8.940 -39.540 ;
        RECT 10.040 -39.590 10.330 -39.540 ;
        RECT 8.650 -39.730 10.330 -39.590 ;
        RECT 8.650 -39.790 8.940 -39.730 ;
        RECT 10.040 -39.790 10.330 -39.730 ;
        RECT 13.370 -39.590 13.660 -39.530 ;
        RECT 14.730 -39.590 15.020 -39.540 ;
        RECT 13.370 -39.730 15.020 -39.590 ;
        RECT 13.370 -39.780 13.660 -39.730 ;
        RECT 14.730 -39.790 15.020 -39.730 ;
        RECT 20.470 -39.590 20.760 -39.540 ;
        RECT 21.860 -39.590 22.150 -39.540 ;
        RECT 20.470 -39.730 22.150 -39.590 ;
        RECT 20.470 -39.790 20.760 -39.730 ;
        RECT 21.860 -39.790 22.150 -39.730 ;
        RECT 25.190 -39.590 25.480 -39.530 ;
        RECT 26.550 -39.590 26.840 -39.540 ;
        RECT 25.190 -39.730 26.840 -39.590 ;
        RECT 25.190 -39.780 25.480 -39.730 ;
        RECT 26.550 -39.790 26.840 -39.730 ;
        RECT 32.290 -39.590 32.580 -39.540 ;
        RECT 33.680 -39.590 33.970 -39.540 ;
        RECT 32.290 -39.730 33.970 -39.590 ;
        RECT 32.290 -39.790 32.580 -39.730 ;
        RECT 33.680 -39.790 33.970 -39.730 ;
        RECT 37.010 -39.590 37.300 -39.530 ;
        RECT 38.370 -39.590 38.660 -39.540 ;
        RECT 37.010 -39.730 38.660 -39.590 ;
        RECT 37.010 -39.780 37.300 -39.730 ;
        RECT 38.370 -39.790 38.660 -39.730 ;
        RECT 44.110 -39.590 44.400 -39.540 ;
        RECT 45.500 -39.590 45.790 -39.540 ;
        RECT 44.110 -39.730 45.790 -39.590 ;
        RECT 44.110 -39.790 44.400 -39.730 ;
        RECT 45.500 -39.790 45.790 -39.730 ;
        RECT 48.830 -39.590 49.120 -39.530 ;
        RECT 50.190 -39.590 50.480 -39.540 ;
        RECT 48.830 -39.730 50.480 -39.590 ;
        RECT 48.830 -39.780 49.120 -39.730 ;
        RECT 50.190 -39.790 50.480 -39.730 ;
        RECT 55.930 -39.590 56.220 -39.540 ;
        RECT 57.320 -39.590 57.610 -39.540 ;
        RECT 55.930 -39.730 57.610 -39.590 ;
        RECT 55.930 -39.790 56.220 -39.730 ;
        RECT 57.320 -39.790 57.610 -39.730 ;
        RECT 60.650 -39.590 60.940 -39.530 ;
        RECT 62.010 -39.590 62.300 -39.540 ;
        RECT 60.650 -39.730 62.300 -39.590 ;
        RECT 60.650 -39.780 60.940 -39.730 ;
        RECT 62.010 -39.790 62.300 -39.730 ;
        RECT 67.750 -39.590 68.040 -39.540 ;
        RECT 69.140 -39.590 69.430 -39.540 ;
        RECT 67.750 -39.730 69.430 -39.590 ;
        RECT 67.750 -39.790 68.040 -39.730 ;
        RECT 69.140 -39.790 69.430 -39.730 ;
        RECT 72.470 -39.590 72.760 -39.530 ;
        RECT 73.830 -39.590 74.120 -39.540 ;
        RECT 72.470 -39.730 74.120 -39.590 ;
        RECT 72.470 -39.780 72.760 -39.730 ;
        RECT 73.830 -39.790 74.120 -39.730 ;
        RECT 79.570 -39.590 79.860 -39.540 ;
        RECT 80.960 -39.590 81.250 -39.540 ;
        RECT 79.570 -39.730 81.250 -39.590 ;
        RECT 79.570 -39.790 79.860 -39.730 ;
        RECT 80.960 -39.790 81.250 -39.730 ;
        RECT 84.290 -39.590 84.580 -39.530 ;
        RECT 85.650 -39.590 85.940 -39.540 ;
        RECT 84.290 -39.730 85.940 -39.590 ;
        RECT 84.290 -39.780 84.580 -39.730 ;
        RECT 85.650 -39.790 85.940 -39.730 ;
        RECT 91.410 -39.590 91.700 -39.540 ;
        RECT 92.800 -39.590 93.090 -39.540 ;
        RECT 91.410 -39.730 93.090 -39.590 ;
        RECT 91.410 -39.790 91.700 -39.730 ;
        RECT 92.800 -39.790 93.090 -39.730 ;
        RECT 96.130 -39.590 96.420 -39.530 ;
        RECT 97.490 -39.590 97.780 -39.540 ;
        RECT 96.130 -39.730 97.780 -39.590 ;
        RECT 96.130 -39.780 96.420 -39.730 ;
        RECT 97.490 -39.790 97.780 -39.730 ;
        RECT 103.250 -39.590 103.540 -39.540 ;
        RECT 104.640 -39.590 104.930 -39.540 ;
        RECT 103.250 -39.730 104.930 -39.590 ;
        RECT 103.250 -39.790 103.540 -39.730 ;
        RECT 104.640 -39.790 104.930 -39.730 ;
        RECT 107.970 -39.590 108.260 -39.530 ;
        RECT 109.330 -39.590 109.620 -39.540 ;
        RECT 107.970 -39.730 109.620 -39.590 ;
        RECT 107.970 -39.780 108.260 -39.730 ;
        RECT 109.330 -39.790 109.620 -39.730 ;
        RECT 115.120 -39.590 115.410 -39.540 ;
        RECT 116.510 -39.590 116.800 -39.540 ;
        RECT 115.120 -39.730 116.800 -39.590 ;
        RECT 115.120 -39.790 115.410 -39.730 ;
        RECT 116.510 -39.790 116.800 -39.730 ;
        RECT 119.840 -39.590 120.130 -39.530 ;
        RECT 121.200 -39.590 121.490 -39.540 ;
        RECT 119.840 -39.730 121.490 -39.590 ;
        RECT 119.840 -39.780 120.130 -39.730 ;
        RECT 121.200 -39.790 121.490 -39.730 ;
        RECT 126.990 -39.590 127.280 -39.540 ;
        RECT 128.380 -39.590 128.670 -39.540 ;
        RECT 126.990 -39.730 128.670 -39.590 ;
        RECT 126.990 -39.790 127.280 -39.730 ;
        RECT 128.380 -39.790 128.670 -39.730 ;
        RECT 131.710 -39.590 132.000 -39.530 ;
        RECT 133.070 -39.590 133.360 -39.540 ;
        RECT 131.710 -39.730 133.360 -39.590 ;
        RECT 131.710 -39.780 132.000 -39.730 ;
        RECT 133.070 -39.790 133.360 -39.730 ;
        RECT 136.000 -39.590 136.290 -39.540 ;
        RECT 137.390 -39.590 137.680 -39.540 ;
        RECT 136.000 -39.730 137.680 -39.590 ;
        RECT 136.000 -39.790 136.290 -39.730 ;
        RECT 137.390 -39.790 137.680 -39.730 ;
        RECT 140.720 -39.590 141.010 -39.530 ;
        RECT 142.080 -39.590 142.370 -39.540 ;
        RECT 140.720 -39.730 142.370 -39.590 ;
        RECT 140.720 -39.780 141.010 -39.730 ;
        RECT 142.080 -39.790 142.370 -39.730 ;
        RECT -39.300 -41.400 -38.920 -41.280 ;
        RECT -37.980 -41.380 -37.680 -41.320 ;
        RECT -37.980 -41.400 -37.670 -41.380 ;
        RECT -39.300 -41.540 -37.670 -41.400 ;
        RECT -39.300 -41.660 -38.920 -41.540 ;
        RECT -37.980 -41.550 -37.670 -41.540 ;
        RECT -27.430 -41.390 -27.170 -41.320 ;
        RECT -26.480 -41.380 -26.180 -41.320 ;
        RECT -27.430 -41.400 -26.940 -41.390 ;
        RECT -26.480 -41.400 -26.170 -41.380 ;
        RECT -27.430 -41.540 -26.170 -41.400 ;
        RECT -37.980 -41.600 -37.680 -41.550 ;
        RECT -27.430 -41.560 -26.940 -41.540 ;
        RECT -26.480 -41.550 -26.170 -41.540 ;
        RECT -15.670 -41.390 -15.350 -41.350 ;
        RECT -14.660 -41.380 -14.360 -41.320 ;
        RECT -15.670 -41.400 -15.120 -41.390 ;
        RECT -14.660 -41.400 -14.350 -41.380 ;
        RECT -15.670 -41.540 -14.350 -41.400 ;
        RECT -27.430 -41.640 -27.170 -41.560 ;
        RECT -26.480 -41.600 -26.180 -41.550 ;
        RECT -15.670 -41.560 -15.120 -41.540 ;
        RECT -14.660 -41.550 -14.350 -41.540 ;
        RECT -3.890 -41.390 -3.570 -41.350 ;
        RECT -2.850 -41.380 -2.550 -41.320 ;
        RECT -3.890 -41.400 -3.310 -41.390 ;
        RECT -2.850 -41.400 -2.540 -41.380 ;
        RECT -3.890 -41.540 -2.540 -41.400 ;
        RECT -15.670 -41.610 -15.350 -41.560 ;
        RECT -14.660 -41.600 -14.360 -41.550 ;
        RECT -3.890 -41.560 -3.310 -41.540 ;
        RECT -2.850 -41.550 -2.540 -41.540 ;
        RECT 8.090 -41.390 8.410 -41.350 ;
        RECT 8.960 -41.380 9.260 -41.320 ;
        RECT 19.760 -41.380 20.080 -41.340 ;
        RECT 20.780 -41.380 21.080 -41.320 ;
        RECT 31.350 -41.370 31.670 -41.330 ;
        RECT 8.090 -41.400 8.500 -41.390 ;
        RECT 8.960 -41.400 9.270 -41.380 ;
        RECT 8.090 -41.540 9.270 -41.400 ;
        RECT -3.890 -41.610 -3.570 -41.560 ;
        RECT -2.850 -41.600 -2.550 -41.550 ;
        RECT 8.090 -41.610 8.410 -41.540 ;
        RECT 8.960 -41.550 9.270 -41.540 ;
        RECT 19.760 -41.400 20.320 -41.380 ;
        RECT 20.780 -41.400 21.090 -41.380 ;
        RECT 19.760 -41.540 21.090 -41.400 ;
        RECT 19.760 -41.550 20.320 -41.540 ;
        RECT 20.780 -41.550 21.090 -41.540 ;
        RECT 31.350 -41.400 32.140 -41.370 ;
        RECT 32.600 -41.380 32.900 -41.320 ;
        RECT 43.090 -41.370 43.410 -41.330 ;
        RECT 32.600 -41.400 32.910 -41.380 ;
        RECT 31.350 -41.540 32.910 -41.400 ;
        RECT 8.960 -41.600 9.260 -41.550 ;
        RECT 19.760 -41.600 20.080 -41.550 ;
        RECT 20.780 -41.600 21.080 -41.550 ;
        RECT 31.350 -41.590 31.670 -41.540 ;
        RECT 32.600 -41.550 32.910 -41.540 ;
        RECT 43.090 -41.400 43.960 -41.370 ;
        RECT 44.420 -41.380 44.720 -41.320 ;
        RECT 54.940 -41.370 55.260 -41.330 ;
        RECT 44.420 -41.400 44.730 -41.380 ;
        RECT 43.090 -41.540 44.730 -41.400 ;
        RECT 32.600 -41.600 32.900 -41.550 ;
        RECT 43.090 -41.590 43.410 -41.540 ;
        RECT 44.420 -41.550 44.730 -41.540 ;
        RECT 54.940 -41.400 55.780 -41.370 ;
        RECT 56.240 -41.380 56.540 -41.320 ;
        RECT 56.240 -41.400 56.550 -41.380 ;
        RECT 54.940 -41.540 56.550 -41.400 ;
        RECT 44.420 -41.600 44.720 -41.550 ;
        RECT 54.940 -41.590 55.260 -41.540 ;
        RECT 56.240 -41.550 56.550 -41.540 ;
        RECT 66.440 -41.390 66.760 -41.350 ;
        RECT 68.060 -41.380 68.360 -41.320 ;
        RECT 66.440 -41.400 67.600 -41.390 ;
        RECT 68.060 -41.400 68.370 -41.380 ;
        RECT 66.440 -41.540 68.370 -41.400 ;
        RECT 56.240 -41.600 56.540 -41.550 ;
        RECT 66.440 -41.560 67.600 -41.540 ;
        RECT 68.060 -41.550 68.370 -41.540 ;
        RECT 78.460 -41.390 78.780 -41.350 ;
        RECT 79.880 -41.380 80.180 -41.320 ;
        RECT 78.460 -41.400 79.420 -41.390 ;
        RECT 79.880 -41.400 80.190 -41.380 ;
        RECT 78.460 -41.540 80.190 -41.400 ;
        RECT 66.440 -41.610 66.760 -41.560 ;
        RECT 68.060 -41.600 68.360 -41.550 ;
        RECT 78.460 -41.560 79.420 -41.540 ;
        RECT 79.880 -41.550 80.190 -41.540 ;
        RECT 90.370 -41.390 90.630 -41.320 ;
        RECT 91.720 -41.380 92.020 -41.320 ;
        RECT 90.370 -41.400 91.260 -41.390 ;
        RECT 91.720 -41.400 92.030 -41.380 ;
        RECT 90.370 -41.540 92.030 -41.400 ;
        RECT 78.460 -41.610 78.780 -41.560 ;
        RECT 79.880 -41.600 80.180 -41.550 ;
        RECT 90.370 -41.560 91.260 -41.540 ;
        RECT 91.720 -41.550 92.030 -41.540 ;
        RECT 102.080 -41.390 102.400 -41.350 ;
        RECT 103.560 -41.380 103.860 -41.320 ;
        RECT 114.210 -41.380 114.530 -41.340 ;
        RECT 115.430 -41.380 115.730 -41.320 ;
        RECT 102.080 -41.400 103.100 -41.390 ;
        RECT 103.560 -41.400 103.870 -41.380 ;
        RECT 102.080 -41.540 103.870 -41.400 ;
        RECT 90.370 -41.640 90.630 -41.560 ;
        RECT 91.720 -41.600 92.020 -41.550 ;
        RECT 102.080 -41.560 103.100 -41.540 ;
        RECT 103.560 -41.550 103.870 -41.540 ;
        RECT 114.210 -41.400 114.970 -41.380 ;
        RECT 115.430 -41.400 115.740 -41.380 ;
        RECT 114.210 -41.540 115.740 -41.400 ;
        RECT 114.210 -41.550 114.970 -41.540 ;
        RECT 115.430 -41.550 115.740 -41.540 ;
        RECT 125.840 -41.390 126.160 -41.350 ;
        RECT 127.300 -41.380 127.600 -41.320 ;
        RECT 135.330 -41.380 135.590 -41.310 ;
        RECT 136.310 -41.380 136.610 -41.320 ;
        RECT 125.840 -41.400 126.840 -41.390 ;
        RECT 127.300 -41.400 127.610 -41.380 ;
        RECT 125.840 -41.540 127.610 -41.400 ;
        RECT 102.080 -41.610 102.400 -41.560 ;
        RECT 103.560 -41.600 103.860 -41.550 ;
        RECT 114.210 -41.600 114.530 -41.550 ;
        RECT 115.430 -41.600 115.730 -41.550 ;
        RECT 125.840 -41.560 126.840 -41.540 ;
        RECT 127.300 -41.550 127.610 -41.540 ;
        RECT 135.330 -41.400 135.850 -41.380 ;
        RECT 136.310 -41.400 136.620 -41.380 ;
        RECT 135.330 -41.540 136.620 -41.400 ;
        RECT 135.330 -41.550 135.850 -41.540 ;
        RECT 136.310 -41.550 136.620 -41.540 ;
        RECT 125.840 -41.610 126.160 -41.560 ;
        RECT 127.300 -41.600 127.600 -41.550 ;
        RECT 135.330 -41.630 135.590 -41.550 ;
        RECT 136.310 -41.600 136.610 -41.550 ;
        RECT -41.810 -43.520 -41.490 -43.460 ;
        RECT -39.160 -43.520 -38.840 -43.460 ;
        RECT -37.490 -43.520 -37.210 -43.450 ;
        RECT -32.940 -43.520 -32.620 -43.460 ;
        RECT -25.990 -43.520 -25.710 -43.450 ;
        RECT -21.440 -43.520 -21.120 -43.460 ;
        RECT -14.170 -43.520 -13.890 -43.450 ;
        RECT -9.620 -43.520 -9.300 -43.460 ;
        RECT -2.360 -43.520 -2.080 -43.450 ;
        RECT 2.190 -43.520 2.510 -43.460 ;
        RECT 9.450 -43.520 9.730 -43.450 ;
        RECT 14.000 -43.520 14.320 -43.460 ;
        RECT 21.270 -43.520 21.550 -43.450 ;
        RECT 25.820 -43.520 26.140 -43.460 ;
        RECT 33.090 -43.520 33.370 -43.450 ;
        RECT 37.640 -43.520 37.960 -43.460 ;
        RECT 44.910 -43.520 45.190 -43.450 ;
        RECT 49.460 -43.520 49.780 -43.460 ;
        RECT 56.730 -43.520 57.010 -43.450 ;
        RECT 61.280 -43.520 61.600 -43.460 ;
        RECT 68.550 -43.520 68.830 -43.450 ;
        RECT 73.100 -43.520 73.420 -43.460 ;
        RECT 80.370 -43.520 80.650 -43.450 ;
        RECT 84.920 -43.520 85.240 -43.460 ;
        RECT 92.210 -43.520 92.490 -43.450 ;
        RECT 96.760 -43.520 97.080 -43.460 ;
        RECT 104.050 -43.520 104.330 -43.450 ;
        RECT 108.600 -43.520 108.920 -43.460 ;
        RECT 115.920 -43.520 116.200 -43.450 ;
        RECT 120.470 -43.520 120.790 -43.460 ;
        RECT 127.790 -43.520 128.070 -43.450 ;
        RECT 132.340 -43.520 132.660 -43.460 ;
        RECT 136.800 -43.520 137.080 -43.450 ;
        RECT 141.350 -43.520 141.670 -43.460 ;
        RECT -41.810 -43.660 142.470 -43.520 ;
        RECT -41.810 -43.720 -41.490 -43.660 ;
        RECT -39.160 -43.720 -38.840 -43.660 ;
        RECT -37.490 -43.750 -37.210 -43.660 ;
        RECT -32.940 -43.720 -32.620 -43.660 ;
        RECT -25.990 -43.750 -25.710 -43.660 ;
        RECT -21.440 -43.720 -21.120 -43.660 ;
        RECT -14.170 -43.750 -13.890 -43.660 ;
        RECT -9.620 -43.720 -9.300 -43.660 ;
        RECT -2.360 -43.750 -2.080 -43.660 ;
        RECT 2.190 -43.720 2.510 -43.660 ;
        RECT 9.450 -43.750 9.730 -43.660 ;
        RECT 14.000 -43.720 14.320 -43.660 ;
        RECT 21.270 -43.750 21.550 -43.660 ;
        RECT 25.820 -43.720 26.140 -43.660 ;
        RECT 33.090 -43.750 33.370 -43.660 ;
        RECT 37.640 -43.720 37.960 -43.660 ;
        RECT 44.910 -43.750 45.190 -43.660 ;
        RECT 49.460 -43.720 49.780 -43.660 ;
        RECT 56.730 -43.750 57.010 -43.660 ;
        RECT 61.280 -43.720 61.600 -43.660 ;
        RECT 68.550 -43.750 68.830 -43.660 ;
        RECT 73.100 -43.720 73.420 -43.660 ;
        RECT 80.370 -43.750 80.650 -43.660 ;
        RECT 84.920 -43.720 85.240 -43.660 ;
        RECT 92.210 -43.750 92.490 -43.660 ;
        RECT 96.760 -43.720 97.080 -43.660 ;
        RECT 104.050 -43.750 104.330 -43.660 ;
        RECT 108.600 -43.720 108.920 -43.660 ;
        RECT 115.920 -43.750 116.200 -43.660 ;
        RECT 120.470 -43.720 120.790 -43.660 ;
        RECT 127.790 -43.750 128.070 -43.660 ;
        RECT 132.340 -43.720 132.660 -43.660 ;
        RECT 136.800 -43.750 137.080 -43.660 ;
        RECT 141.350 -43.720 141.670 -43.660 ;
        RECT -37.860 -43.920 -37.620 -43.910 ;
        RECT -26.360 -43.920 -26.120 -43.910 ;
        RECT -14.540 -43.920 -14.300 -43.910 ;
        RECT -2.730 -43.920 -2.490 -43.910 ;
        RECT 9.080 -43.920 9.320 -43.910 ;
        RECT 20.900 -43.920 21.140 -43.910 ;
        RECT 32.720 -43.920 32.960 -43.910 ;
        RECT 44.540 -43.920 44.780 -43.910 ;
        RECT 56.360 -43.920 56.600 -43.910 ;
        RECT 68.180 -43.920 68.420 -43.910 ;
        RECT 80.000 -43.920 80.240 -43.910 ;
        RECT 91.840 -43.920 92.080 -43.910 ;
        RECT 103.680 -43.920 103.920 -43.910 ;
        RECT 115.550 -43.920 115.790 -43.910 ;
        RECT 127.420 -43.920 127.660 -43.910 ;
        RECT 136.430 -43.920 136.670 -43.910 ;
        RECT -37.900 -44.240 -37.580 -43.920 ;
        RECT -26.400 -44.240 -26.080 -43.920 ;
        RECT -14.580 -44.240 -14.260 -43.920 ;
        RECT -2.770 -44.240 -2.450 -43.920 ;
        RECT 9.040 -44.240 9.360 -43.920 ;
        RECT 20.860 -44.240 21.180 -43.920 ;
        RECT 32.680 -44.240 33.000 -43.920 ;
        RECT 44.500 -44.240 44.820 -43.920 ;
        RECT 56.320 -44.240 56.640 -43.920 ;
        RECT 68.140 -44.240 68.460 -43.920 ;
        RECT 79.960 -44.240 80.280 -43.920 ;
        RECT 91.800 -44.240 92.120 -43.920 ;
        RECT 103.640 -44.240 103.960 -43.920 ;
        RECT 115.510 -44.240 115.830 -43.920 ;
        RECT 127.380 -44.240 127.700 -43.920 ;
        RECT 136.390 -44.240 136.710 -43.920 ;
        RECT -32.210 -44.500 -31.920 -44.480 ;
        RECT -20.710 -44.500 -20.420 -44.470 ;
        RECT -8.890 -44.500 -8.600 -44.470 ;
        RECT 2.920 -44.500 3.210 -44.470 ;
        RECT 14.730 -44.500 15.020 -44.470 ;
        RECT 26.550 -44.500 26.840 -44.470 ;
        RECT 38.370 -44.500 38.660 -44.470 ;
        RECT 50.190 -44.500 50.480 -44.470 ;
        RECT 62.010 -44.500 62.300 -44.470 ;
        RECT 73.830 -44.500 74.120 -44.470 ;
        RECT 85.650 -44.500 85.940 -44.470 ;
        RECT 97.490 -44.500 97.780 -44.470 ;
        RECT 109.330 -44.500 109.620 -44.470 ;
        RECT 121.200 -44.500 121.490 -44.470 ;
        RECT 133.070 -44.500 133.360 -44.470 ;
        RECT 142.110 -44.500 142.340 -44.440 ;
        RECT 144.430 -44.500 144.750 -44.450 ;
        RECT -32.210 -44.670 144.750 -44.500 ;
        RECT -32.210 -44.710 -31.920 -44.670 ;
        RECT -20.710 -44.700 -20.420 -44.670 ;
        RECT -8.890 -44.700 -8.600 -44.670 ;
        RECT 2.920 -44.700 3.210 -44.670 ;
        RECT 14.730 -44.700 15.020 -44.670 ;
        RECT 26.550 -44.700 26.840 -44.670 ;
        RECT 38.370 -44.700 38.660 -44.670 ;
        RECT 50.190 -44.700 50.480 -44.670 ;
        RECT 62.010 -44.700 62.300 -44.670 ;
        RECT 73.830 -44.700 74.120 -44.670 ;
        RECT 85.650 -44.700 85.940 -44.670 ;
        RECT 97.490 -44.700 97.780 -44.670 ;
        RECT 109.330 -44.700 109.620 -44.670 ;
        RECT 121.200 -44.700 121.490 -44.670 ;
        RECT 133.070 -44.700 133.360 -44.670 ;
        RECT 142.110 -44.730 142.340 -44.670 ;
        RECT 144.430 -44.710 144.750 -44.670 ;
        RECT -32.940 -45.230 -32.580 -44.890 ;
        RECT -21.440 -45.230 -21.080 -44.890 ;
        RECT -9.620 -45.230 -9.260 -44.890 ;
        RECT 2.190 -45.230 2.550 -44.890 ;
        RECT 14.000 -45.230 14.360 -44.890 ;
        RECT 25.820 -45.230 26.180 -44.890 ;
        RECT 37.640 -45.230 38.000 -44.890 ;
        RECT 49.460 -45.230 49.820 -44.890 ;
        RECT 61.280 -45.230 61.640 -44.890 ;
        RECT 73.100 -45.230 73.460 -44.890 ;
        RECT 84.920 -45.230 85.280 -44.890 ;
        RECT 96.760 -45.230 97.120 -44.890 ;
        RECT 108.600 -45.230 108.960 -44.890 ;
        RECT 120.470 -45.230 120.830 -44.890 ;
        RECT 132.340 -45.230 132.700 -44.890 ;
        RECT 141.350 -45.230 141.710 -44.890 ;
        RECT -32.210 -45.390 -31.920 -45.370 ;
        RECT -20.710 -45.390 -20.420 -45.360 ;
        RECT 2.920 -45.390 3.210 -45.360 ;
        RECT 14.730 -45.390 15.020 -45.360 ;
        RECT 26.550 -45.390 26.840 -45.360 ;
        RECT 38.370 -45.390 38.660 -45.360 ;
        RECT 50.190 -45.390 50.480 -45.360 ;
        RECT 62.010 -45.390 62.300 -45.360 ;
        RECT 73.830 -45.390 74.120 -45.360 ;
        RECT 85.650 -45.390 85.940 -45.360 ;
        RECT 97.490 -45.390 97.780 -45.360 ;
        RECT 109.330 -45.390 109.620 -45.370 ;
        RECT 121.200 -45.390 121.490 -45.360 ;
        RECT 133.070 -45.390 133.360 -45.360 ;
        RECT 142.080 -45.390 142.370 -45.360 ;
        RECT 144.990 -45.390 145.310 -45.340 ;
        RECT -32.210 -45.560 145.310 -45.390 ;
        RECT -32.210 -45.600 -31.920 -45.560 ;
        RECT -20.710 -45.590 -20.420 -45.560 ;
        RECT -8.890 -45.620 -8.600 -45.560 ;
        RECT 2.920 -45.590 3.210 -45.560 ;
        RECT 14.730 -45.590 15.020 -45.560 ;
        RECT 26.550 -45.590 26.840 -45.560 ;
        RECT 38.370 -45.590 38.660 -45.560 ;
        RECT 50.190 -45.590 50.480 -45.560 ;
        RECT 62.010 -45.590 62.300 -45.560 ;
        RECT 73.830 -45.590 74.120 -45.560 ;
        RECT 85.650 -45.590 85.940 -45.560 ;
        RECT 97.490 -45.590 97.780 -45.560 ;
        RECT 109.330 -45.600 109.620 -45.560 ;
        RECT 121.200 -45.590 121.490 -45.560 ;
        RECT 133.070 -45.590 133.360 -45.560 ;
        RECT 142.080 -45.590 142.370 -45.560 ;
        RECT 144.990 -45.600 145.310 -45.560 ;
        RECT -39.160 -46.420 -38.840 -46.360 ;
        RECT -37.490 -46.420 -37.210 -46.330 ;
        RECT -32.910 -46.420 -32.650 -46.330 ;
        RECT -25.990 -46.420 -25.710 -46.330 ;
        RECT -21.410 -46.420 -21.150 -46.330 ;
        RECT -14.170 -46.420 -13.890 -46.330 ;
        RECT -9.590 -46.420 -9.330 -46.330 ;
        RECT -2.360 -46.420 -2.080 -46.330 ;
        RECT 2.220 -46.420 2.480 -46.330 ;
        RECT 9.450 -46.420 9.730 -46.330 ;
        RECT 14.030 -46.420 14.290 -46.330 ;
        RECT 21.270 -46.420 21.550 -46.330 ;
        RECT 25.850 -46.420 26.110 -46.330 ;
        RECT 33.090 -46.420 33.370 -46.330 ;
        RECT 37.670 -46.420 37.930 -46.330 ;
        RECT 44.910 -46.420 45.190 -46.330 ;
        RECT 49.490 -46.420 49.750 -46.330 ;
        RECT 56.730 -46.420 57.010 -46.330 ;
        RECT 61.310 -46.420 61.570 -46.330 ;
        RECT 68.550 -46.420 68.830 -46.330 ;
        RECT 73.130 -46.420 73.390 -46.330 ;
        RECT 80.370 -46.420 80.650 -46.330 ;
        RECT 84.950 -46.420 85.210 -46.330 ;
        RECT 92.210 -46.420 92.490 -46.330 ;
        RECT 96.790 -46.420 97.050 -46.330 ;
        RECT 104.050 -46.420 104.330 -46.330 ;
        RECT 108.630 -46.420 108.890 -46.330 ;
        RECT 115.920 -46.420 116.200 -46.330 ;
        RECT 120.500 -46.420 120.760 -46.330 ;
        RECT 127.790 -46.420 128.070 -46.330 ;
        RECT 132.370 -46.420 132.630 -46.330 ;
        RECT 136.800 -46.420 137.080 -46.330 ;
        RECT 141.380 -46.420 141.640 -46.330 ;
        RECT -39.160 -46.560 142.470 -46.420 ;
        RECT -39.160 -46.620 -38.840 -46.560 ;
        RECT -37.490 -46.630 -37.210 -46.560 ;
        RECT -32.910 -46.650 -32.650 -46.560 ;
        RECT -25.990 -46.630 -25.710 -46.560 ;
        RECT -21.410 -46.650 -21.150 -46.560 ;
        RECT -14.170 -46.630 -13.890 -46.560 ;
        RECT -9.590 -46.650 -9.330 -46.560 ;
        RECT -2.360 -46.630 -2.080 -46.560 ;
        RECT 2.220 -46.650 2.480 -46.560 ;
        RECT 9.450 -46.630 9.730 -46.560 ;
        RECT 14.030 -46.650 14.290 -46.560 ;
        RECT 21.270 -46.630 21.550 -46.560 ;
        RECT 25.850 -46.650 26.110 -46.560 ;
        RECT 33.090 -46.630 33.370 -46.560 ;
        RECT 37.670 -46.650 37.930 -46.560 ;
        RECT 44.910 -46.630 45.190 -46.560 ;
        RECT 49.490 -46.650 49.750 -46.560 ;
        RECT 56.730 -46.630 57.010 -46.560 ;
        RECT 61.310 -46.650 61.570 -46.560 ;
        RECT 68.550 -46.630 68.830 -46.560 ;
        RECT 73.130 -46.650 73.390 -46.560 ;
        RECT 80.370 -46.630 80.650 -46.560 ;
        RECT 84.950 -46.650 85.210 -46.560 ;
        RECT 92.210 -46.630 92.490 -46.560 ;
        RECT 96.790 -46.650 97.050 -46.560 ;
        RECT 104.050 -46.630 104.330 -46.560 ;
        RECT 108.630 -46.650 108.890 -46.560 ;
        RECT 115.920 -46.630 116.200 -46.560 ;
        RECT 120.500 -46.650 120.760 -46.560 ;
        RECT 127.790 -46.630 128.070 -46.560 ;
        RECT 132.370 -46.650 132.630 -46.560 ;
        RECT 136.800 -46.630 137.080 -46.560 ;
        RECT 141.380 -46.650 141.640 -46.560 ;
        RECT -37.910 -48.780 -37.590 -48.460 ;
        RECT -26.410 -48.780 -26.090 -48.460 ;
        RECT -14.590 -48.780 -14.270 -48.460 ;
        RECT -2.780 -48.780 -2.460 -48.460 ;
        RECT 9.030 -48.780 9.350 -48.460 ;
        RECT 20.850 -48.780 21.170 -48.460 ;
        RECT 32.670 -48.780 32.990 -48.460 ;
        RECT 44.490 -48.780 44.810 -48.460 ;
        RECT 56.310 -48.780 56.630 -48.460 ;
        RECT 68.130 -48.780 68.450 -48.460 ;
        RECT 79.950 -48.780 80.270 -48.460 ;
        RECT 91.790 -48.780 92.110 -48.460 ;
        RECT 103.630 -48.780 103.950 -48.460 ;
        RECT 115.500 -48.780 115.820 -48.460 ;
        RECT 127.370 -48.780 127.690 -48.460 ;
        RECT 136.380 -48.780 136.700 -48.460 ;
        RECT -37.870 -48.790 -37.630 -48.780 ;
        RECT -26.370 -48.790 -26.130 -48.780 ;
        RECT -14.550 -48.790 -14.310 -48.780 ;
        RECT -2.740 -48.790 -2.500 -48.780 ;
        RECT 9.070 -48.790 9.310 -48.780 ;
        RECT 20.890 -48.790 21.130 -48.780 ;
        RECT 32.710 -48.790 32.950 -48.780 ;
        RECT 44.530 -48.790 44.770 -48.780 ;
        RECT 56.350 -48.790 56.590 -48.780 ;
        RECT 68.170 -48.790 68.410 -48.780 ;
        RECT 79.990 -48.790 80.230 -48.780 ;
        RECT 91.830 -48.790 92.070 -48.780 ;
        RECT 103.670 -48.790 103.910 -48.780 ;
        RECT 115.540 -48.790 115.780 -48.780 ;
        RECT 127.410 -48.790 127.650 -48.780 ;
        RECT 136.420 -48.790 136.660 -48.780 ;
        RECT -38.290 -50.350 -38.000 -50.290 ;
        RECT -36.900 -50.350 -36.610 -50.290 ;
        RECT -38.290 -50.490 -36.610 -50.350 ;
        RECT -38.290 -50.540 -38.000 -50.490 ;
        RECT -36.900 -50.540 -36.610 -50.490 ;
        RECT -33.570 -50.350 -33.280 -50.300 ;
        RECT -32.210 -50.350 -31.920 -50.290 ;
        RECT -33.570 -50.490 -31.920 -50.350 ;
        RECT -33.570 -50.550 -33.280 -50.490 ;
        RECT -32.210 -50.540 -31.920 -50.490 ;
        RECT -26.790 -50.350 -26.500 -50.290 ;
        RECT -25.400 -50.350 -25.110 -50.290 ;
        RECT -26.790 -50.490 -25.110 -50.350 ;
        RECT -26.790 -50.540 -26.500 -50.490 ;
        RECT -25.400 -50.540 -25.110 -50.490 ;
        RECT -22.070 -50.350 -21.780 -50.300 ;
        RECT -20.710 -50.350 -20.420 -50.290 ;
        RECT -22.070 -50.490 -20.420 -50.350 ;
        RECT -22.070 -50.550 -21.780 -50.490 ;
        RECT -20.710 -50.540 -20.420 -50.490 ;
        RECT -14.970 -50.350 -14.680 -50.290 ;
        RECT -13.580 -50.350 -13.290 -50.290 ;
        RECT -14.970 -50.490 -13.290 -50.350 ;
        RECT -14.970 -50.540 -14.680 -50.490 ;
        RECT -13.580 -50.540 -13.290 -50.490 ;
        RECT -10.250 -50.350 -9.960 -50.300 ;
        RECT -8.890 -50.350 -8.600 -50.290 ;
        RECT -10.250 -50.490 -8.600 -50.350 ;
        RECT -10.250 -50.550 -9.960 -50.490 ;
        RECT -8.890 -50.540 -8.600 -50.490 ;
        RECT -3.160 -50.350 -2.870 -50.290 ;
        RECT -1.770 -50.350 -1.480 -50.290 ;
        RECT -3.160 -50.490 -1.480 -50.350 ;
        RECT -3.160 -50.540 -2.870 -50.490 ;
        RECT -1.770 -50.540 -1.480 -50.490 ;
        RECT 1.560 -50.350 1.850 -50.300 ;
        RECT 2.920 -50.350 3.210 -50.290 ;
        RECT 1.560 -50.490 3.210 -50.350 ;
        RECT 1.560 -50.550 1.850 -50.490 ;
        RECT 2.920 -50.540 3.210 -50.490 ;
        RECT 8.650 -50.350 8.940 -50.290 ;
        RECT 10.040 -50.350 10.330 -50.290 ;
        RECT 8.650 -50.490 10.330 -50.350 ;
        RECT 8.650 -50.540 8.940 -50.490 ;
        RECT 10.040 -50.540 10.330 -50.490 ;
        RECT 13.370 -50.350 13.660 -50.300 ;
        RECT 14.730 -50.350 15.020 -50.290 ;
        RECT 13.370 -50.490 15.020 -50.350 ;
        RECT 13.370 -50.550 13.660 -50.490 ;
        RECT 14.730 -50.540 15.020 -50.490 ;
        RECT 20.470 -50.350 20.760 -50.290 ;
        RECT 21.860 -50.350 22.150 -50.290 ;
        RECT 20.470 -50.490 22.150 -50.350 ;
        RECT 20.470 -50.540 20.760 -50.490 ;
        RECT 21.860 -50.540 22.150 -50.490 ;
        RECT 25.190 -50.350 25.480 -50.300 ;
        RECT 26.550 -50.350 26.840 -50.290 ;
        RECT 25.190 -50.490 26.840 -50.350 ;
        RECT 25.190 -50.550 25.480 -50.490 ;
        RECT 26.550 -50.540 26.840 -50.490 ;
        RECT 32.290 -50.350 32.580 -50.290 ;
        RECT 33.680 -50.350 33.970 -50.290 ;
        RECT 32.290 -50.490 33.970 -50.350 ;
        RECT 32.290 -50.540 32.580 -50.490 ;
        RECT 33.680 -50.540 33.970 -50.490 ;
        RECT 37.010 -50.350 37.300 -50.300 ;
        RECT 38.370 -50.350 38.660 -50.290 ;
        RECT 37.010 -50.490 38.660 -50.350 ;
        RECT 37.010 -50.550 37.300 -50.490 ;
        RECT 38.370 -50.540 38.660 -50.490 ;
        RECT 44.110 -50.350 44.400 -50.290 ;
        RECT 45.500 -50.350 45.790 -50.290 ;
        RECT 44.110 -50.490 45.790 -50.350 ;
        RECT 44.110 -50.540 44.400 -50.490 ;
        RECT 45.500 -50.540 45.790 -50.490 ;
        RECT 48.830 -50.350 49.120 -50.300 ;
        RECT 50.190 -50.350 50.480 -50.290 ;
        RECT 48.830 -50.490 50.480 -50.350 ;
        RECT 48.830 -50.550 49.120 -50.490 ;
        RECT 50.190 -50.540 50.480 -50.490 ;
        RECT 55.930 -50.350 56.220 -50.290 ;
        RECT 57.320 -50.350 57.610 -50.290 ;
        RECT 55.930 -50.490 57.610 -50.350 ;
        RECT 55.930 -50.540 56.220 -50.490 ;
        RECT 57.320 -50.540 57.610 -50.490 ;
        RECT 60.650 -50.350 60.940 -50.300 ;
        RECT 62.010 -50.350 62.300 -50.290 ;
        RECT 60.650 -50.490 62.300 -50.350 ;
        RECT 60.650 -50.550 60.940 -50.490 ;
        RECT 62.010 -50.540 62.300 -50.490 ;
        RECT 67.750 -50.350 68.040 -50.290 ;
        RECT 69.140 -50.350 69.430 -50.290 ;
        RECT 67.750 -50.490 69.430 -50.350 ;
        RECT 67.750 -50.540 68.040 -50.490 ;
        RECT 69.140 -50.540 69.430 -50.490 ;
        RECT 72.470 -50.350 72.760 -50.300 ;
        RECT 73.830 -50.350 74.120 -50.290 ;
        RECT 72.470 -50.490 74.120 -50.350 ;
        RECT 72.470 -50.550 72.760 -50.490 ;
        RECT 73.830 -50.540 74.120 -50.490 ;
        RECT 79.570 -50.350 79.860 -50.290 ;
        RECT 80.960 -50.350 81.250 -50.290 ;
        RECT 79.570 -50.490 81.250 -50.350 ;
        RECT 79.570 -50.540 79.860 -50.490 ;
        RECT 80.960 -50.540 81.250 -50.490 ;
        RECT 84.290 -50.350 84.580 -50.300 ;
        RECT 85.650 -50.350 85.940 -50.290 ;
        RECT 84.290 -50.490 85.940 -50.350 ;
        RECT 84.290 -50.550 84.580 -50.490 ;
        RECT 85.650 -50.540 85.940 -50.490 ;
        RECT 91.410 -50.350 91.700 -50.290 ;
        RECT 92.800 -50.350 93.090 -50.290 ;
        RECT 91.410 -50.490 93.090 -50.350 ;
        RECT 91.410 -50.540 91.700 -50.490 ;
        RECT 92.800 -50.540 93.090 -50.490 ;
        RECT 96.130 -50.350 96.420 -50.300 ;
        RECT 97.490 -50.350 97.780 -50.290 ;
        RECT 96.130 -50.490 97.780 -50.350 ;
        RECT 96.130 -50.550 96.420 -50.490 ;
        RECT 97.490 -50.540 97.780 -50.490 ;
        RECT 103.250 -50.350 103.540 -50.290 ;
        RECT 104.640 -50.350 104.930 -50.290 ;
        RECT 103.250 -50.490 104.930 -50.350 ;
        RECT 103.250 -50.540 103.540 -50.490 ;
        RECT 104.640 -50.540 104.930 -50.490 ;
        RECT 107.970 -50.350 108.260 -50.300 ;
        RECT 109.330 -50.350 109.620 -50.290 ;
        RECT 107.970 -50.490 109.620 -50.350 ;
        RECT 107.970 -50.550 108.260 -50.490 ;
        RECT 109.330 -50.540 109.620 -50.490 ;
        RECT 115.120 -50.350 115.410 -50.290 ;
        RECT 116.510 -50.350 116.800 -50.290 ;
        RECT 115.120 -50.490 116.800 -50.350 ;
        RECT 115.120 -50.540 115.410 -50.490 ;
        RECT 116.510 -50.540 116.800 -50.490 ;
        RECT 119.840 -50.350 120.130 -50.300 ;
        RECT 121.200 -50.350 121.490 -50.290 ;
        RECT 119.840 -50.490 121.490 -50.350 ;
        RECT 119.840 -50.550 120.130 -50.490 ;
        RECT 121.200 -50.540 121.490 -50.490 ;
        RECT 126.990 -50.350 127.280 -50.290 ;
        RECT 128.380 -50.350 128.670 -50.290 ;
        RECT 126.990 -50.490 128.670 -50.350 ;
        RECT 126.990 -50.540 127.280 -50.490 ;
        RECT 128.380 -50.540 128.670 -50.490 ;
        RECT 131.710 -50.350 132.000 -50.300 ;
        RECT 133.070 -50.350 133.360 -50.290 ;
        RECT 131.710 -50.490 133.360 -50.350 ;
        RECT 131.710 -50.550 132.000 -50.490 ;
        RECT 133.070 -50.540 133.360 -50.490 ;
        RECT 136.000 -50.350 136.290 -50.290 ;
        RECT 137.390 -50.350 137.680 -50.290 ;
        RECT 136.000 -50.490 137.680 -50.350 ;
        RECT 136.000 -50.540 136.290 -50.490 ;
        RECT 137.390 -50.540 137.680 -50.490 ;
        RECT 140.720 -50.350 141.010 -50.300 ;
        RECT 142.080 -50.350 142.370 -50.290 ;
        RECT 140.720 -50.490 142.370 -50.350 ;
        RECT 140.720 -50.550 141.010 -50.490 ;
        RECT 142.080 -50.540 142.370 -50.490 ;
        RECT -34.970 -51.090 -34.680 -51.030 ;
        RECT -34.010 -51.090 -33.720 -51.020 ;
        RECT -34.970 -51.230 -33.720 -51.090 ;
        RECT -34.970 -51.280 -34.680 -51.230 ;
        RECT -34.010 -51.270 -33.720 -51.230 ;
        RECT -23.470 -51.090 -23.180 -51.030 ;
        RECT -22.510 -51.090 -22.220 -51.020 ;
        RECT -23.470 -51.230 -22.220 -51.090 ;
        RECT -23.470 -51.280 -23.180 -51.230 ;
        RECT -22.510 -51.270 -22.220 -51.230 ;
        RECT -11.650 -51.090 -11.360 -51.030 ;
        RECT -10.690 -51.090 -10.400 -51.020 ;
        RECT -11.650 -51.230 -10.400 -51.090 ;
        RECT -11.650 -51.280 -11.360 -51.230 ;
        RECT -10.690 -51.270 -10.400 -51.230 ;
        RECT 0.160 -51.090 0.450 -51.030 ;
        RECT 1.120 -51.090 1.410 -51.020 ;
        RECT 0.160 -51.230 1.410 -51.090 ;
        RECT 0.160 -51.280 0.450 -51.230 ;
        RECT 1.120 -51.270 1.410 -51.230 ;
        RECT 11.970 -51.090 12.260 -51.030 ;
        RECT 12.930 -51.090 13.220 -51.020 ;
        RECT 11.970 -51.230 13.220 -51.090 ;
        RECT 11.970 -51.280 12.260 -51.230 ;
        RECT 12.930 -51.270 13.220 -51.230 ;
        RECT 23.790 -51.090 24.080 -51.030 ;
        RECT 24.750 -51.090 25.040 -51.020 ;
        RECT 23.790 -51.230 25.040 -51.090 ;
        RECT 23.790 -51.280 24.080 -51.230 ;
        RECT 24.750 -51.270 25.040 -51.230 ;
        RECT 35.610 -51.090 35.900 -51.030 ;
        RECT 36.570 -51.090 36.860 -51.020 ;
        RECT 35.610 -51.230 36.860 -51.090 ;
        RECT 35.610 -51.280 35.900 -51.230 ;
        RECT 36.570 -51.270 36.860 -51.230 ;
        RECT 47.430 -51.090 47.720 -51.030 ;
        RECT 48.390 -51.090 48.680 -51.020 ;
        RECT 47.430 -51.230 48.680 -51.090 ;
        RECT 47.430 -51.280 47.720 -51.230 ;
        RECT 48.390 -51.270 48.680 -51.230 ;
        RECT 59.250 -51.090 59.540 -51.030 ;
        RECT 60.210 -51.090 60.500 -51.020 ;
        RECT 59.250 -51.230 60.500 -51.090 ;
        RECT 59.250 -51.280 59.540 -51.230 ;
        RECT 60.210 -51.270 60.500 -51.230 ;
        RECT 71.070 -51.090 71.360 -51.030 ;
        RECT 72.030 -51.090 72.320 -51.020 ;
        RECT 71.070 -51.230 72.320 -51.090 ;
        RECT 71.070 -51.280 71.360 -51.230 ;
        RECT 72.030 -51.270 72.320 -51.230 ;
        RECT 82.890 -51.090 83.180 -51.030 ;
        RECT 83.850 -51.090 84.140 -51.020 ;
        RECT 82.890 -51.230 84.140 -51.090 ;
        RECT 82.890 -51.280 83.180 -51.230 ;
        RECT 83.850 -51.270 84.140 -51.230 ;
        RECT 94.730 -51.090 95.020 -51.030 ;
        RECT 95.690 -51.090 95.980 -51.020 ;
        RECT 94.730 -51.230 95.980 -51.090 ;
        RECT 94.730 -51.280 95.020 -51.230 ;
        RECT 95.690 -51.270 95.980 -51.230 ;
        RECT 106.570 -51.090 106.860 -51.030 ;
        RECT 107.530 -51.090 107.820 -51.020 ;
        RECT 106.570 -51.230 107.820 -51.090 ;
        RECT 106.570 -51.280 106.860 -51.230 ;
        RECT 107.530 -51.270 107.820 -51.230 ;
        RECT 118.440 -51.090 118.730 -51.030 ;
        RECT 119.400 -51.090 119.690 -51.020 ;
        RECT 118.440 -51.230 119.690 -51.090 ;
        RECT 118.440 -51.280 118.730 -51.230 ;
        RECT 119.400 -51.270 119.690 -51.230 ;
        RECT 130.310 -51.090 130.600 -51.030 ;
        RECT 131.270 -51.090 131.560 -51.020 ;
        RECT 130.310 -51.230 131.560 -51.090 ;
        RECT 130.310 -51.280 130.600 -51.230 ;
        RECT 131.270 -51.270 131.560 -51.230 ;
        RECT 139.320 -51.090 139.610 -51.030 ;
        RECT 140.280 -51.090 140.570 -51.020 ;
        RECT 139.320 -51.230 140.570 -51.090 ;
        RECT 139.320 -51.280 139.610 -51.230 ;
        RECT 140.280 -51.270 140.570 -51.230 ;
        RECT -36.460 -51.900 -36.170 -51.840 ;
        RECT -35.500 -51.900 -35.210 -51.840 ;
        RECT -36.460 -52.040 -35.210 -51.900 ;
        RECT -36.460 -52.090 -36.170 -52.040 ;
        RECT -35.500 -52.090 -35.210 -52.040 ;
        RECT -24.960 -51.900 -24.670 -51.840 ;
        RECT -24.000 -51.900 -23.710 -51.840 ;
        RECT -24.960 -52.040 -23.710 -51.900 ;
        RECT -24.960 -52.090 -24.670 -52.040 ;
        RECT -24.000 -52.090 -23.710 -52.040 ;
        RECT -13.140 -51.900 -12.850 -51.840 ;
        RECT -12.180 -51.900 -11.890 -51.840 ;
        RECT -13.140 -52.040 -11.890 -51.900 ;
        RECT -13.140 -52.090 -12.850 -52.040 ;
        RECT -12.180 -52.090 -11.890 -52.040 ;
        RECT -1.330 -51.900 -1.040 -51.840 ;
        RECT -0.370 -51.900 -0.080 -51.840 ;
        RECT -1.330 -52.040 -0.080 -51.900 ;
        RECT -1.330 -52.090 -1.040 -52.040 ;
        RECT -0.370 -52.090 -0.080 -52.040 ;
        RECT 10.480 -51.900 10.770 -51.840 ;
        RECT 11.440 -51.900 11.730 -51.840 ;
        RECT 10.480 -52.040 11.730 -51.900 ;
        RECT 10.480 -52.090 10.770 -52.040 ;
        RECT 11.440 -52.090 11.730 -52.040 ;
        RECT 22.300 -51.900 22.590 -51.840 ;
        RECT 23.260 -51.900 23.550 -51.840 ;
        RECT 22.300 -52.040 23.550 -51.900 ;
        RECT 22.300 -52.090 22.590 -52.040 ;
        RECT 23.260 -52.090 23.550 -52.040 ;
        RECT 34.120 -51.900 34.410 -51.840 ;
        RECT 35.080 -51.900 35.370 -51.840 ;
        RECT 34.120 -52.040 35.370 -51.900 ;
        RECT 34.120 -52.090 34.410 -52.040 ;
        RECT 35.080 -52.090 35.370 -52.040 ;
        RECT 45.940 -51.900 46.230 -51.840 ;
        RECT 46.900 -51.900 47.190 -51.840 ;
        RECT 45.940 -52.040 47.190 -51.900 ;
        RECT 45.940 -52.090 46.230 -52.040 ;
        RECT 46.900 -52.090 47.190 -52.040 ;
        RECT 57.760 -51.900 58.050 -51.840 ;
        RECT 58.720 -51.900 59.010 -51.840 ;
        RECT 57.760 -52.040 59.010 -51.900 ;
        RECT 57.760 -52.090 58.050 -52.040 ;
        RECT 58.720 -52.090 59.010 -52.040 ;
        RECT 69.580 -51.900 69.870 -51.840 ;
        RECT 70.540 -51.900 70.830 -51.840 ;
        RECT 69.580 -52.040 70.830 -51.900 ;
        RECT 69.580 -52.090 69.870 -52.040 ;
        RECT 70.540 -52.090 70.830 -52.040 ;
        RECT 81.400 -51.900 81.690 -51.840 ;
        RECT 82.360 -51.900 82.650 -51.840 ;
        RECT 81.400 -52.040 82.650 -51.900 ;
        RECT 81.400 -52.090 81.690 -52.040 ;
        RECT 82.360 -52.090 82.650 -52.040 ;
        RECT 93.240 -51.900 93.530 -51.840 ;
        RECT 94.200 -51.900 94.490 -51.840 ;
        RECT 93.240 -52.040 94.490 -51.900 ;
        RECT 93.240 -52.090 93.530 -52.040 ;
        RECT 94.200 -52.090 94.490 -52.040 ;
        RECT 105.080 -51.900 105.370 -51.840 ;
        RECT 106.040 -51.900 106.330 -51.840 ;
        RECT 105.080 -52.040 106.330 -51.900 ;
        RECT 105.080 -52.090 105.370 -52.040 ;
        RECT 106.040 -52.090 106.330 -52.040 ;
        RECT 116.950 -51.900 117.240 -51.840 ;
        RECT 117.910 -51.900 118.200 -51.840 ;
        RECT 116.950 -52.040 118.200 -51.900 ;
        RECT 116.950 -52.090 117.240 -52.040 ;
        RECT 117.910 -52.090 118.200 -52.040 ;
        RECT 128.820 -51.900 129.110 -51.840 ;
        RECT 129.780 -51.900 130.070 -51.840 ;
        RECT 128.820 -52.040 130.070 -51.900 ;
        RECT 128.820 -52.090 129.110 -52.040 ;
        RECT 129.780 -52.090 130.070 -52.040 ;
        RECT 137.830 -51.900 138.120 -51.840 ;
        RECT 138.790 -51.900 139.080 -51.840 ;
        RECT 137.830 -52.040 139.080 -51.900 ;
        RECT 137.830 -52.090 138.120 -52.040 ;
        RECT 138.790 -52.090 139.080 -52.040 ;
        RECT -37.940 -52.570 -37.650 -52.520 ;
        RECT -36.460 -52.570 -36.170 -52.550 ;
        RECT -37.940 -52.710 -36.170 -52.570 ;
        RECT -37.940 -52.770 -37.650 -52.710 ;
        RECT -36.460 -52.800 -36.170 -52.710 ;
        RECT -34.010 -52.600 -33.720 -52.560 ;
        RECT -32.560 -52.600 -32.270 -52.530 ;
        RECT -34.010 -52.740 -32.270 -52.600 ;
        RECT -34.010 -52.810 -33.720 -52.740 ;
        RECT -32.560 -52.780 -32.270 -52.740 ;
        RECT -26.440 -52.570 -26.150 -52.520 ;
        RECT -24.960 -52.570 -24.670 -52.550 ;
        RECT -26.440 -52.710 -24.670 -52.570 ;
        RECT -26.440 -52.770 -26.150 -52.710 ;
        RECT -24.960 -52.800 -24.670 -52.710 ;
        RECT -22.510 -52.600 -22.220 -52.560 ;
        RECT -21.060 -52.600 -20.770 -52.530 ;
        RECT -22.510 -52.740 -20.770 -52.600 ;
        RECT -22.510 -52.810 -22.220 -52.740 ;
        RECT -21.060 -52.780 -20.770 -52.740 ;
        RECT -14.620 -52.570 -14.330 -52.520 ;
        RECT -13.140 -52.570 -12.850 -52.550 ;
        RECT -14.620 -52.710 -12.850 -52.570 ;
        RECT -14.620 -52.770 -14.330 -52.710 ;
        RECT -13.140 -52.800 -12.850 -52.710 ;
        RECT -10.690 -52.600 -10.400 -52.560 ;
        RECT -9.240 -52.600 -8.950 -52.530 ;
        RECT -10.690 -52.740 -8.950 -52.600 ;
        RECT -10.690 -52.810 -10.400 -52.740 ;
        RECT -9.240 -52.780 -8.950 -52.740 ;
        RECT -2.810 -52.570 -2.520 -52.520 ;
        RECT -1.330 -52.570 -1.040 -52.550 ;
        RECT -2.810 -52.710 -1.040 -52.570 ;
        RECT -2.810 -52.770 -2.520 -52.710 ;
        RECT -1.330 -52.800 -1.040 -52.710 ;
        RECT 1.120 -52.600 1.410 -52.560 ;
        RECT 2.570 -52.600 2.860 -52.530 ;
        RECT 1.120 -52.740 2.860 -52.600 ;
        RECT 1.120 -52.810 1.410 -52.740 ;
        RECT 2.570 -52.780 2.860 -52.740 ;
        RECT 9.000 -52.570 9.290 -52.520 ;
        RECT 10.480 -52.570 10.770 -52.550 ;
        RECT 9.000 -52.710 10.770 -52.570 ;
        RECT 9.000 -52.770 9.290 -52.710 ;
        RECT 10.480 -52.800 10.770 -52.710 ;
        RECT 12.930 -52.600 13.220 -52.560 ;
        RECT 14.380 -52.600 14.670 -52.530 ;
        RECT 12.930 -52.740 14.670 -52.600 ;
        RECT 12.930 -52.810 13.220 -52.740 ;
        RECT 14.380 -52.780 14.670 -52.740 ;
        RECT 20.820 -52.570 21.110 -52.520 ;
        RECT 22.300 -52.570 22.590 -52.550 ;
        RECT 20.820 -52.710 22.590 -52.570 ;
        RECT 20.820 -52.770 21.110 -52.710 ;
        RECT 22.300 -52.800 22.590 -52.710 ;
        RECT 24.750 -52.600 25.040 -52.560 ;
        RECT 26.200 -52.600 26.490 -52.530 ;
        RECT 24.750 -52.740 26.490 -52.600 ;
        RECT 24.750 -52.810 25.040 -52.740 ;
        RECT 26.200 -52.780 26.490 -52.740 ;
        RECT 32.640 -52.570 32.930 -52.520 ;
        RECT 34.120 -52.570 34.410 -52.550 ;
        RECT 32.640 -52.710 34.410 -52.570 ;
        RECT 32.640 -52.770 32.930 -52.710 ;
        RECT 34.120 -52.800 34.410 -52.710 ;
        RECT 36.570 -52.600 36.860 -52.560 ;
        RECT 38.020 -52.600 38.310 -52.530 ;
        RECT 36.570 -52.740 38.310 -52.600 ;
        RECT 36.570 -52.810 36.860 -52.740 ;
        RECT 38.020 -52.780 38.310 -52.740 ;
        RECT 44.460 -52.570 44.750 -52.520 ;
        RECT 45.940 -52.570 46.230 -52.550 ;
        RECT 44.460 -52.710 46.230 -52.570 ;
        RECT 44.460 -52.770 44.750 -52.710 ;
        RECT 45.940 -52.800 46.230 -52.710 ;
        RECT 48.390 -52.600 48.680 -52.560 ;
        RECT 49.840 -52.600 50.130 -52.530 ;
        RECT 48.390 -52.740 50.130 -52.600 ;
        RECT 48.390 -52.810 48.680 -52.740 ;
        RECT 49.840 -52.780 50.130 -52.740 ;
        RECT 56.280 -52.570 56.570 -52.520 ;
        RECT 57.760 -52.570 58.050 -52.550 ;
        RECT 56.280 -52.710 58.050 -52.570 ;
        RECT 56.280 -52.770 56.570 -52.710 ;
        RECT 57.760 -52.800 58.050 -52.710 ;
        RECT 60.210 -52.600 60.500 -52.560 ;
        RECT 61.660 -52.600 61.950 -52.530 ;
        RECT 60.210 -52.740 61.950 -52.600 ;
        RECT 60.210 -52.810 60.500 -52.740 ;
        RECT 61.660 -52.780 61.950 -52.740 ;
        RECT 68.100 -52.570 68.390 -52.520 ;
        RECT 69.580 -52.570 69.870 -52.550 ;
        RECT 68.100 -52.710 69.870 -52.570 ;
        RECT 68.100 -52.770 68.390 -52.710 ;
        RECT 69.580 -52.800 69.870 -52.710 ;
        RECT 72.030 -52.600 72.320 -52.560 ;
        RECT 73.480 -52.600 73.770 -52.530 ;
        RECT 72.030 -52.740 73.770 -52.600 ;
        RECT 72.030 -52.810 72.320 -52.740 ;
        RECT 73.480 -52.780 73.770 -52.740 ;
        RECT 79.920 -52.570 80.210 -52.520 ;
        RECT 81.400 -52.570 81.690 -52.550 ;
        RECT 79.920 -52.710 81.690 -52.570 ;
        RECT 79.920 -52.770 80.210 -52.710 ;
        RECT 81.400 -52.800 81.690 -52.710 ;
        RECT 83.850 -52.600 84.140 -52.560 ;
        RECT 85.300 -52.600 85.590 -52.530 ;
        RECT 83.850 -52.740 85.590 -52.600 ;
        RECT 83.850 -52.810 84.140 -52.740 ;
        RECT 85.300 -52.780 85.590 -52.740 ;
        RECT 91.760 -52.570 92.050 -52.520 ;
        RECT 93.240 -52.570 93.530 -52.550 ;
        RECT 91.760 -52.710 93.530 -52.570 ;
        RECT 91.760 -52.770 92.050 -52.710 ;
        RECT 93.240 -52.800 93.530 -52.710 ;
        RECT 95.690 -52.600 95.980 -52.560 ;
        RECT 97.140 -52.600 97.430 -52.530 ;
        RECT 95.690 -52.740 97.430 -52.600 ;
        RECT 95.690 -52.810 95.980 -52.740 ;
        RECT 97.140 -52.780 97.430 -52.740 ;
        RECT 103.600 -52.570 103.890 -52.520 ;
        RECT 105.080 -52.570 105.370 -52.550 ;
        RECT 103.600 -52.710 105.370 -52.570 ;
        RECT 103.600 -52.770 103.890 -52.710 ;
        RECT 105.080 -52.800 105.370 -52.710 ;
        RECT 107.530 -52.600 107.820 -52.560 ;
        RECT 108.980 -52.600 109.270 -52.530 ;
        RECT 107.530 -52.740 109.270 -52.600 ;
        RECT 107.530 -52.810 107.820 -52.740 ;
        RECT 108.980 -52.780 109.270 -52.740 ;
        RECT 115.470 -52.570 115.760 -52.520 ;
        RECT 116.950 -52.570 117.240 -52.550 ;
        RECT 115.470 -52.710 117.240 -52.570 ;
        RECT 115.470 -52.770 115.760 -52.710 ;
        RECT 116.950 -52.800 117.240 -52.710 ;
        RECT 119.400 -52.600 119.690 -52.560 ;
        RECT 120.850 -52.600 121.140 -52.530 ;
        RECT 119.400 -52.740 121.140 -52.600 ;
        RECT 119.400 -52.810 119.690 -52.740 ;
        RECT 120.850 -52.780 121.140 -52.740 ;
        RECT 127.340 -52.570 127.630 -52.520 ;
        RECT 128.820 -52.570 129.110 -52.550 ;
        RECT 127.340 -52.710 129.110 -52.570 ;
        RECT 127.340 -52.770 127.630 -52.710 ;
        RECT 128.820 -52.800 129.110 -52.710 ;
        RECT 131.270 -52.600 131.560 -52.560 ;
        RECT 132.720 -52.600 133.010 -52.530 ;
        RECT 131.270 -52.740 133.010 -52.600 ;
        RECT 131.270 -52.810 131.560 -52.740 ;
        RECT 132.720 -52.780 133.010 -52.740 ;
        RECT 136.350 -52.570 136.640 -52.520 ;
        RECT 137.830 -52.570 138.120 -52.550 ;
        RECT 136.350 -52.710 138.120 -52.570 ;
        RECT 136.350 -52.770 136.640 -52.710 ;
        RECT 137.830 -52.800 138.120 -52.710 ;
        RECT 140.280 -52.600 140.570 -52.560 ;
        RECT 141.730 -52.600 142.020 -52.530 ;
        RECT 140.280 -52.740 142.020 -52.600 ;
        RECT 140.280 -52.810 140.570 -52.740 ;
        RECT 141.730 -52.780 142.020 -52.740 ;
        RECT -41.230 -53.200 -40.910 -53.140 ;
        RECT -37.860 -53.190 -37.570 -53.160 ;
        RECT -37.900 -53.200 -37.570 -53.190 ;
        RECT -32.640 -53.170 -32.350 -53.140 ;
        RECT -32.640 -53.200 -32.310 -53.170 ;
        RECT -26.360 -53.190 -26.070 -53.160 ;
        RECT -26.400 -53.200 -26.070 -53.190 ;
        RECT -21.140 -53.170 -20.850 -53.140 ;
        RECT -21.140 -53.200 -20.810 -53.170 ;
        RECT -14.540 -53.190 -14.250 -53.160 ;
        RECT -14.580 -53.200 -14.250 -53.190 ;
        RECT -9.320 -53.170 -9.030 -53.140 ;
        RECT -9.320 -53.200 -8.990 -53.170 ;
        RECT -2.730 -53.190 -2.440 -53.160 ;
        RECT -2.770 -53.200 -2.440 -53.190 ;
        RECT 2.490 -53.170 2.780 -53.140 ;
        RECT 2.490 -53.200 2.820 -53.170 ;
        RECT 9.080 -53.190 9.370 -53.160 ;
        RECT 9.040 -53.200 9.370 -53.190 ;
        RECT 14.300 -53.170 14.590 -53.140 ;
        RECT 14.300 -53.200 14.630 -53.170 ;
        RECT 20.900 -53.190 21.190 -53.160 ;
        RECT 20.860 -53.200 21.190 -53.190 ;
        RECT 26.120 -53.170 26.410 -53.140 ;
        RECT 26.120 -53.200 26.450 -53.170 ;
        RECT 32.720 -53.190 33.010 -53.160 ;
        RECT 32.680 -53.200 33.010 -53.190 ;
        RECT 37.940 -53.170 38.230 -53.140 ;
        RECT 37.940 -53.200 38.270 -53.170 ;
        RECT 44.540 -53.190 44.830 -53.160 ;
        RECT 44.500 -53.200 44.830 -53.190 ;
        RECT 49.760 -53.170 50.050 -53.140 ;
        RECT 49.760 -53.200 50.090 -53.170 ;
        RECT 56.360 -53.190 56.650 -53.160 ;
        RECT 56.320 -53.200 56.650 -53.190 ;
        RECT 61.580 -53.170 61.870 -53.140 ;
        RECT 61.580 -53.200 61.910 -53.170 ;
        RECT 68.180 -53.190 68.470 -53.160 ;
        RECT 68.140 -53.200 68.470 -53.190 ;
        RECT 73.400 -53.170 73.690 -53.140 ;
        RECT 73.400 -53.200 73.730 -53.170 ;
        RECT 80.000 -53.190 80.290 -53.160 ;
        RECT 79.960 -53.200 80.290 -53.190 ;
        RECT 85.220 -53.170 85.510 -53.140 ;
        RECT 85.220 -53.200 85.550 -53.170 ;
        RECT 91.840 -53.190 92.130 -53.160 ;
        RECT 91.800 -53.200 92.130 -53.190 ;
        RECT 97.060 -53.170 97.350 -53.140 ;
        RECT 97.060 -53.200 97.390 -53.170 ;
        RECT 103.680 -53.190 103.970 -53.160 ;
        RECT 103.640 -53.200 103.970 -53.190 ;
        RECT 108.900 -53.170 109.190 -53.140 ;
        RECT 108.900 -53.200 109.230 -53.170 ;
        RECT 115.550 -53.190 115.840 -53.160 ;
        RECT 115.510 -53.200 115.840 -53.190 ;
        RECT 120.770 -53.170 121.060 -53.140 ;
        RECT 120.770 -53.200 121.100 -53.170 ;
        RECT 127.420 -53.190 127.710 -53.160 ;
        RECT 127.380 -53.200 127.710 -53.190 ;
        RECT 132.640 -53.170 132.930 -53.140 ;
        RECT 132.640 -53.200 132.970 -53.170 ;
        RECT 136.430 -53.190 136.720 -53.160 ;
        RECT 136.390 -53.200 136.720 -53.190 ;
        RECT 141.650 -53.170 141.940 -53.140 ;
        RECT 141.650 -53.200 141.980 -53.170 ;
        RECT -41.230 -53.340 142.470 -53.200 ;
        RECT -41.230 -53.400 -40.910 -53.340 ;
        RECT -37.900 -53.370 -37.570 -53.340 ;
        RECT -37.860 -53.400 -37.570 -53.370 ;
        RECT -32.640 -53.350 -32.310 -53.340 ;
        RECT -32.640 -53.380 -32.350 -53.350 ;
        RECT -26.400 -53.370 -26.070 -53.340 ;
        RECT -26.360 -53.400 -26.070 -53.370 ;
        RECT -21.140 -53.350 -20.810 -53.340 ;
        RECT -21.140 -53.380 -20.850 -53.350 ;
        RECT -14.580 -53.370 -14.250 -53.340 ;
        RECT -14.540 -53.400 -14.250 -53.370 ;
        RECT -9.320 -53.350 -8.990 -53.340 ;
        RECT -9.320 -53.380 -9.030 -53.350 ;
        RECT -2.770 -53.370 -2.440 -53.340 ;
        RECT -2.730 -53.400 -2.440 -53.370 ;
        RECT 2.490 -53.350 2.820 -53.340 ;
        RECT 2.490 -53.380 2.780 -53.350 ;
        RECT 9.040 -53.370 9.370 -53.340 ;
        RECT 9.080 -53.400 9.370 -53.370 ;
        RECT 14.300 -53.350 14.630 -53.340 ;
        RECT 14.300 -53.380 14.590 -53.350 ;
        RECT 20.860 -53.370 21.190 -53.340 ;
        RECT 20.900 -53.400 21.190 -53.370 ;
        RECT 26.120 -53.350 26.450 -53.340 ;
        RECT 26.120 -53.380 26.410 -53.350 ;
        RECT 32.680 -53.370 33.010 -53.340 ;
        RECT 32.720 -53.400 33.010 -53.370 ;
        RECT 37.940 -53.350 38.270 -53.340 ;
        RECT 37.940 -53.380 38.230 -53.350 ;
        RECT 44.500 -53.370 44.830 -53.340 ;
        RECT 44.540 -53.400 44.830 -53.370 ;
        RECT 49.760 -53.350 50.090 -53.340 ;
        RECT 49.760 -53.380 50.050 -53.350 ;
        RECT 56.320 -53.370 56.650 -53.340 ;
        RECT 56.360 -53.400 56.650 -53.370 ;
        RECT 61.580 -53.350 61.910 -53.340 ;
        RECT 61.580 -53.380 61.870 -53.350 ;
        RECT 68.140 -53.370 68.470 -53.340 ;
        RECT 68.180 -53.400 68.470 -53.370 ;
        RECT 73.400 -53.350 73.730 -53.340 ;
        RECT 73.400 -53.380 73.690 -53.350 ;
        RECT 79.960 -53.370 80.290 -53.340 ;
        RECT 80.000 -53.400 80.290 -53.370 ;
        RECT 85.220 -53.350 85.550 -53.340 ;
        RECT 85.220 -53.380 85.510 -53.350 ;
        RECT 91.800 -53.370 92.130 -53.340 ;
        RECT 91.840 -53.400 92.130 -53.370 ;
        RECT 97.060 -53.350 97.390 -53.340 ;
        RECT 97.060 -53.380 97.350 -53.350 ;
        RECT 103.640 -53.370 103.970 -53.340 ;
        RECT 103.680 -53.400 103.970 -53.370 ;
        RECT 108.900 -53.350 109.230 -53.340 ;
        RECT 108.900 -53.380 109.190 -53.350 ;
        RECT 115.510 -53.370 115.840 -53.340 ;
        RECT 115.550 -53.400 115.840 -53.370 ;
        RECT 120.770 -53.350 121.100 -53.340 ;
        RECT 120.770 -53.380 121.060 -53.350 ;
        RECT 127.380 -53.370 127.710 -53.340 ;
        RECT 127.420 -53.400 127.710 -53.370 ;
        RECT 132.640 -53.350 132.970 -53.340 ;
        RECT 132.640 -53.380 132.930 -53.350 ;
        RECT 136.390 -53.370 136.720 -53.340 ;
        RECT 136.430 -53.400 136.720 -53.370 ;
        RECT 141.650 -53.350 141.980 -53.340 ;
        RECT 141.650 -53.380 141.940 -53.350 ;
        RECT -40.570 -53.600 -40.250 -53.540 ;
        RECT -36.790 -53.600 -36.460 -53.550 ;
        RECT -33.720 -53.600 -33.390 -53.560 ;
        RECT -25.290 -53.600 -24.960 -53.550 ;
        RECT -22.220 -53.600 -21.890 -53.560 ;
        RECT -13.470 -53.600 -13.140 -53.550 ;
        RECT -10.400 -53.600 -10.070 -53.560 ;
        RECT -1.660 -53.600 -1.330 -53.550 ;
        RECT 1.410 -53.600 1.740 -53.560 ;
        RECT 10.150 -53.600 10.480 -53.550 ;
        RECT 13.220 -53.600 13.550 -53.560 ;
        RECT 21.970 -53.600 22.300 -53.550 ;
        RECT 25.040 -53.600 25.370 -53.560 ;
        RECT 33.790 -53.600 34.120 -53.550 ;
        RECT 36.860 -53.600 37.190 -53.560 ;
        RECT 45.610 -53.600 45.940 -53.550 ;
        RECT 48.680 -53.600 49.010 -53.560 ;
        RECT 57.430 -53.600 57.760 -53.550 ;
        RECT 60.500 -53.600 60.830 -53.560 ;
        RECT 69.250 -53.600 69.580 -53.550 ;
        RECT 72.320 -53.600 72.650 -53.560 ;
        RECT 81.070 -53.600 81.400 -53.550 ;
        RECT 84.140 -53.600 84.470 -53.560 ;
        RECT 92.910 -53.600 93.240 -53.550 ;
        RECT 95.980 -53.600 96.310 -53.560 ;
        RECT 104.750 -53.600 105.080 -53.550 ;
        RECT 107.820 -53.600 108.150 -53.560 ;
        RECT 116.620 -53.600 116.950 -53.550 ;
        RECT 119.690 -53.600 120.020 -53.560 ;
        RECT 128.490 -53.600 128.820 -53.550 ;
        RECT 131.560 -53.600 131.890 -53.560 ;
        RECT 137.500 -53.600 137.830 -53.550 ;
        RECT 140.570 -53.600 140.900 -53.560 ;
        RECT -40.570 -53.740 142.470 -53.600 ;
        RECT -40.570 -53.800 -40.250 -53.740 ;
        RECT -36.790 -53.790 -36.460 -53.740 ;
        RECT -33.720 -53.800 -33.390 -53.740 ;
        RECT -25.290 -53.790 -24.960 -53.740 ;
        RECT -22.220 -53.800 -21.890 -53.740 ;
        RECT -13.470 -53.790 -13.140 -53.740 ;
        RECT -10.400 -53.800 -10.070 -53.740 ;
        RECT -1.660 -53.790 -1.330 -53.740 ;
        RECT 1.410 -53.800 1.740 -53.740 ;
        RECT 10.150 -53.790 10.480 -53.740 ;
        RECT 13.220 -53.800 13.550 -53.740 ;
        RECT 21.970 -53.790 22.300 -53.740 ;
        RECT 25.040 -53.800 25.370 -53.740 ;
        RECT 33.790 -53.790 34.120 -53.740 ;
        RECT 36.860 -53.800 37.190 -53.740 ;
        RECT 45.610 -53.790 45.940 -53.740 ;
        RECT 48.680 -53.800 49.010 -53.740 ;
        RECT 57.430 -53.790 57.760 -53.740 ;
        RECT 60.500 -53.800 60.830 -53.740 ;
        RECT 69.250 -53.790 69.580 -53.740 ;
        RECT 72.320 -53.800 72.650 -53.740 ;
        RECT 81.070 -53.790 81.400 -53.740 ;
        RECT 84.140 -53.800 84.470 -53.740 ;
        RECT 92.910 -53.790 93.240 -53.740 ;
        RECT 95.980 -53.800 96.310 -53.740 ;
        RECT 104.750 -53.790 105.080 -53.740 ;
        RECT 107.820 -53.800 108.150 -53.740 ;
        RECT 116.620 -53.790 116.950 -53.740 ;
        RECT 119.690 -53.800 120.020 -53.740 ;
        RECT 128.490 -53.790 128.820 -53.740 ;
        RECT 131.560 -53.800 131.890 -53.740 ;
        RECT 137.500 -53.790 137.830 -53.740 ;
        RECT 140.570 -53.800 140.900 -53.740 ;
        RECT -36.380 -54.030 -36.090 -53.980 ;
        RECT -31.100 -54.030 -30.780 -53.970 ;
        RECT -36.380 -54.170 -30.780 -54.030 ;
        RECT -36.380 -54.210 -36.090 -54.170 ;
        RECT -31.100 -54.230 -30.780 -54.170 ;
        RECT -25.070 -54.030 -24.780 -53.960 ;
        RECT -19.560 -54.030 -19.240 -53.970 ;
        RECT -25.070 -54.170 -19.240 -54.030 ;
        RECT -25.070 -54.250 -24.780 -54.170 ;
        RECT -19.560 -54.230 -19.240 -54.170 ;
        RECT -13.260 -54.030 -12.970 -53.960 ;
        RECT -7.870 -54.030 -7.550 -53.970 ;
        RECT -13.260 -54.170 -7.550 -54.030 ;
        RECT -13.260 -54.250 -12.970 -54.170 ;
        RECT -7.870 -54.230 -7.550 -54.170 ;
        RECT -1.540 -54.030 -1.250 -53.960 ;
        RECT 4.040 -54.030 4.360 -53.970 ;
        RECT -1.540 -54.170 4.360 -54.030 ;
        RECT -1.540 -54.250 -1.250 -54.170 ;
        RECT 4.040 -54.230 4.360 -54.170 ;
        RECT 10.240 -54.030 10.530 -53.960 ;
        RECT 15.810 -54.030 16.130 -53.970 ;
        RECT 10.240 -54.170 16.130 -54.030 ;
        RECT 10.240 -54.250 10.530 -54.170 ;
        RECT 15.810 -54.230 16.130 -54.170 ;
        RECT 22.120 -54.030 22.410 -53.960 ;
        RECT 27.580 -54.030 27.900 -53.970 ;
        RECT 22.120 -54.170 27.900 -54.030 ;
        RECT 22.120 -54.250 22.410 -54.170 ;
        RECT 27.580 -54.230 27.900 -54.170 ;
        RECT 34.030 -54.030 34.320 -53.960 ;
        RECT 39.400 -54.030 39.720 -53.970 ;
        RECT 34.030 -54.170 39.720 -54.030 ;
        RECT 34.030 -54.250 34.320 -54.170 ;
        RECT 39.400 -54.230 39.720 -54.170 ;
        RECT 45.880 -54.030 46.110 -53.960 ;
        RECT 51.260 -54.030 51.580 -53.970 ;
        RECT 45.880 -54.170 51.580 -54.030 ;
        RECT 45.880 -54.250 46.110 -54.170 ;
        RECT 51.260 -54.230 51.580 -54.170 ;
        RECT 57.540 -54.030 57.830 -53.960 ;
        RECT 63.050 -54.030 63.370 -53.970 ;
        RECT 57.540 -54.170 63.370 -54.030 ;
        RECT 57.540 -54.250 57.830 -54.170 ;
        RECT 63.050 -54.230 63.370 -54.170 ;
        RECT 69.420 -54.030 69.710 -53.960 ;
        RECT 74.930 -54.030 75.250 -53.970 ;
        RECT 69.420 -54.170 75.250 -54.030 ;
        RECT 69.420 -54.250 69.710 -54.170 ;
        RECT 74.930 -54.230 75.250 -54.170 ;
        RECT 81.210 -54.030 81.500 -53.960 ;
        RECT 86.660 -54.030 86.980 -53.970 ;
        RECT 81.210 -54.170 86.980 -54.030 ;
        RECT 81.210 -54.250 81.500 -54.170 ;
        RECT 86.660 -54.230 86.980 -54.170 ;
        RECT 93.090 -54.030 93.380 -53.960 ;
        RECT 98.480 -54.030 98.800 -53.970 ;
        RECT 93.090 -54.170 98.800 -54.030 ;
        RECT 93.090 -54.250 93.380 -54.170 ;
        RECT 98.480 -54.230 98.800 -54.170 ;
        RECT 104.860 -54.030 105.150 -53.960 ;
        RECT 110.370 -54.030 110.690 -53.970 ;
        RECT 104.860 -54.170 110.690 -54.030 ;
        RECT 104.860 -54.250 105.150 -54.170 ;
        RECT 110.370 -54.230 110.690 -54.170 ;
        RECT 116.640 -54.030 116.930 -53.960 ;
        RECT 122.320 -54.030 122.640 -53.970 ;
        RECT 116.640 -54.170 122.640 -54.030 ;
        RECT 116.640 -54.250 116.930 -54.170 ;
        RECT 122.320 -54.230 122.640 -54.170 ;
        RECT 128.450 -54.030 128.740 -53.960 ;
        RECT 134.080 -54.030 134.400 -53.970 ;
        RECT 128.450 -54.170 134.400 -54.030 ;
        RECT 128.450 -54.250 128.740 -54.170 ;
        RECT 134.080 -54.230 134.400 -54.170 ;
        RECT 137.720 -54.030 138.010 -53.960 ;
        RECT 143.120 -54.030 143.440 -53.970 ;
        RECT 137.720 -54.170 143.440 -54.030 ;
        RECT 137.720 -54.250 138.010 -54.170 ;
        RECT 143.120 -54.230 143.440 -54.170 ;
        RECT -37.000 -56.270 -36.750 -56.160 ;
        RECT -35.250 -56.270 -34.930 -56.180 ;
        RECT -37.000 -56.280 -34.930 -56.270 ;
        RECT -33.460 -56.280 -33.210 -56.190 ;
        RECT -32.350 -56.280 -32.060 -56.230 ;
        RECT -37.000 -56.410 -32.060 -56.280 ;
        RECT -37.000 -56.520 -36.750 -56.410 ;
        RECT -35.250 -56.420 -32.060 -56.410 ;
        RECT -35.250 -56.500 -34.930 -56.420 ;
        RECT -33.460 -56.510 -33.210 -56.420 ;
        RECT -32.350 -56.460 -32.060 -56.420 ;
        RECT -25.500 -56.270 -25.250 -56.160 ;
        RECT -23.750 -56.270 -23.430 -56.180 ;
        RECT -25.500 -56.280 -23.430 -56.270 ;
        RECT -21.960 -56.280 -21.710 -56.190 ;
        RECT -20.850 -56.280 -20.560 -56.230 ;
        RECT -25.500 -56.410 -20.560 -56.280 ;
        RECT -25.500 -56.520 -25.250 -56.410 ;
        RECT -23.750 -56.420 -20.560 -56.410 ;
        RECT -23.750 -56.500 -23.430 -56.420 ;
        RECT -21.960 -56.510 -21.710 -56.420 ;
        RECT -20.850 -56.460 -20.560 -56.420 ;
        RECT -13.680 -56.270 -13.430 -56.160 ;
        RECT -11.930 -56.270 -11.610 -56.180 ;
        RECT -13.680 -56.280 -11.610 -56.270 ;
        RECT -10.140 -56.280 -9.890 -56.190 ;
        RECT -9.030 -56.280 -8.740 -56.230 ;
        RECT -13.680 -56.410 -8.740 -56.280 ;
        RECT -13.680 -56.520 -13.430 -56.410 ;
        RECT -11.930 -56.420 -8.740 -56.410 ;
        RECT -11.930 -56.500 -11.610 -56.420 ;
        RECT -10.140 -56.510 -9.890 -56.420 ;
        RECT -9.030 -56.460 -8.740 -56.420 ;
        RECT -1.870 -56.270 -1.620 -56.160 ;
        RECT -0.120 -56.270 0.200 -56.180 ;
        RECT -1.870 -56.280 0.200 -56.270 ;
        RECT 1.670 -56.280 1.920 -56.190 ;
        RECT 2.780 -56.280 3.070 -56.230 ;
        RECT -1.870 -56.410 3.070 -56.280 ;
        RECT -1.870 -56.520 -1.620 -56.410 ;
        RECT -0.120 -56.420 3.070 -56.410 ;
        RECT -0.120 -56.500 0.200 -56.420 ;
        RECT 1.670 -56.510 1.920 -56.420 ;
        RECT 2.780 -56.460 3.070 -56.420 ;
        RECT 9.940 -56.270 10.190 -56.160 ;
        RECT 11.690 -56.270 12.010 -56.180 ;
        RECT 9.940 -56.280 12.010 -56.270 ;
        RECT 13.480 -56.280 13.730 -56.190 ;
        RECT 14.590 -56.280 14.880 -56.230 ;
        RECT 9.940 -56.410 14.880 -56.280 ;
        RECT 9.940 -56.520 10.190 -56.410 ;
        RECT 11.690 -56.420 14.880 -56.410 ;
        RECT 11.690 -56.500 12.010 -56.420 ;
        RECT 13.480 -56.510 13.730 -56.420 ;
        RECT 14.590 -56.460 14.880 -56.420 ;
        RECT 21.760 -56.270 22.010 -56.160 ;
        RECT 23.510 -56.270 23.830 -56.180 ;
        RECT 21.760 -56.280 23.830 -56.270 ;
        RECT 25.300 -56.280 25.550 -56.190 ;
        RECT 26.410 -56.280 26.700 -56.230 ;
        RECT 21.760 -56.410 26.700 -56.280 ;
        RECT 21.760 -56.520 22.010 -56.410 ;
        RECT 23.510 -56.420 26.700 -56.410 ;
        RECT 23.510 -56.500 23.830 -56.420 ;
        RECT 25.300 -56.510 25.550 -56.420 ;
        RECT 26.410 -56.460 26.700 -56.420 ;
        RECT 33.580 -56.270 33.830 -56.160 ;
        RECT 35.330 -56.270 35.650 -56.180 ;
        RECT 33.580 -56.280 35.650 -56.270 ;
        RECT 37.120 -56.280 37.370 -56.190 ;
        RECT 38.230 -56.280 38.520 -56.230 ;
        RECT 33.580 -56.410 38.520 -56.280 ;
        RECT 33.580 -56.520 33.830 -56.410 ;
        RECT 35.330 -56.420 38.520 -56.410 ;
        RECT 35.330 -56.500 35.650 -56.420 ;
        RECT 37.120 -56.510 37.370 -56.420 ;
        RECT 38.230 -56.460 38.520 -56.420 ;
        RECT 45.400 -56.270 45.650 -56.160 ;
        RECT 47.150 -56.270 47.470 -56.180 ;
        RECT 45.400 -56.280 47.470 -56.270 ;
        RECT 48.940 -56.280 49.190 -56.190 ;
        RECT 50.050 -56.280 50.340 -56.230 ;
        RECT 45.400 -56.410 50.340 -56.280 ;
        RECT 45.400 -56.520 45.650 -56.410 ;
        RECT 47.150 -56.420 50.340 -56.410 ;
        RECT 47.150 -56.500 47.470 -56.420 ;
        RECT 48.940 -56.510 49.190 -56.420 ;
        RECT 50.050 -56.460 50.340 -56.420 ;
        RECT 57.220 -56.270 57.470 -56.160 ;
        RECT 58.970 -56.270 59.290 -56.180 ;
        RECT 57.220 -56.280 59.290 -56.270 ;
        RECT 60.760 -56.280 61.010 -56.190 ;
        RECT 61.870 -56.280 62.160 -56.230 ;
        RECT 57.220 -56.410 62.160 -56.280 ;
        RECT 57.220 -56.520 57.470 -56.410 ;
        RECT 58.970 -56.420 62.160 -56.410 ;
        RECT 58.970 -56.500 59.290 -56.420 ;
        RECT 60.760 -56.510 61.010 -56.420 ;
        RECT 61.870 -56.460 62.160 -56.420 ;
        RECT 69.040 -56.270 69.290 -56.160 ;
        RECT 70.790 -56.270 71.110 -56.180 ;
        RECT 69.040 -56.280 71.110 -56.270 ;
        RECT 72.580 -56.280 72.830 -56.190 ;
        RECT 73.690 -56.280 73.980 -56.230 ;
        RECT 69.040 -56.410 73.980 -56.280 ;
        RECT 69.040 -56.520 69.290 -56.410 ;
        RECT 70.790 -56.420 73.980 -56.410 ;
        RECT 70.790 -56.500 71.110 -56.420 ;
        RECT 72.580 -56.510 72.830 -56.420 ;
        RECT 73.690 -56.460 73.980 -56.420 ;
        RECT 80.860 -56.270 81.110 -56.160 ;
        RECT 82.610 -56.270 82.930 -56.180 ;
        RECT 80.860 -56.280 82.930 -56.270 ;
        RECT 84.400 -56.280 84.650 -56.190 ;
        RECT 85.510 -56.280 85.800 -56.230 ;
        RECT 80.860 -56.410 85.800 -56.280 ;
        RECT 80.860 -56.520 81.110 -56.410 ;
        RECT 82.610 -56.420 85.800 -56.410 ;
        RECT 82.610 -56.500 82.930 -56.420 ;
        RECT 84.400 -56.510 84.650 -56.420 ;
        RECT 85.510 -56.460 85.800 -56.420 ;
        RECT 92.700 -56.270 92.950 -56.160 ;
        RECT 94.450 -56.270 94.770 -56.180 ;
        RECT 92.700 -56.280 94.770 -56.270 ;
        RECT 96.240 -56.280 96.490 -56.190 ;
        RECT 97.350 -56.280 97.640 -56.230 ;
        RECT 92.700 -56.410 97.640 -56.280 ;
        RECT 92.700 -56.520 92.950 -56.410 ;
        RECT 94.450 -56.420 97.640 -56.410 ;
        RECT 94.450 -56.500 94.770 -56.420 ;
        RECT 96.240 -56.510 96.490 -56.420 ;
        RECT 97.350 -56.460 97.640 -56.420 ;
        RECT 104.540 -56.270 104.790 -56.160 ;
        RECT 106.290 -56.270 106.610 -56.180 ;
        RECT 104.540 -56.280 106.610 -56.270 ;
        RECT 108.080 -56.280 108.330 -56.190 ;
        RECT 109.190 -56.280 109.480 -56.230 ;
        RECT 104.540 -56.410 109.480 -56.280 ;
        RECT 104.540 -56.520 104.790 -56.410 ;
        RECT 106.290 -56.420 109.480 -56.410 ;
        RECT 106.290 -56.500 106.610 -56.420 ;
        RECT 108.080 -56.510 108.330 -56.420 ;
        RECT 109.190 -56.460 109.480 -56.420 ;
        RECT 116.410 -56.270 116.660 -56.160 ;
        RECT 118.160 -56.270 118.480 -56.180 ;
        RECT 116.410 -56.280 118.480 -56.270 ;
        RECT 119.950 -56.280 120.200 -56.190 ;
        RECT 121.060 -56.280 121.350 -56.230 ;
        RECT 116.410 -56.410 121.350 -56.280 ;
        RECT 116.410 -56.520 116.660 -56.410 ;
        RECT 118.160 -56.420 121.350 -56.410 ;
        RECT 118.160 -56.500 118.480 -56.420 ;
        RECT 119.950 -56.510 120.200 -56.420 ;
        RECT 121.060 -56.460 121.350 -56.420 ;
        RECT 128.280 -56.270 128.530 -56.160 ;
        RECT 130.030 -56.270 130.350 -56.180 ;
        RECT 128.280 -56.280 130.350 -56.270 ;
        RECT 131.820 -56.280 132.070 -56.190 ;
        RECT 132.930 -56.280 133.220 -56.230 ;
        RECT 128.280 -56.410 133.220 -56.280 ;
        RECT 128.280 -56.520 128.530 -56.410 ;
        RECT 130.030 -56.420 133.220 -56.410 ;
        RECT 130.030 -56.500 130.350 -56.420 ;
        RECT 131.820 -56.510 132.070 -56.420 ;
        RECT 132.930 -56.460 133.220 -56.420 ;
        RECT 137.290 -56.270 137.540 -56.160 ;
        RECT 139.040 -56.270 139.360 -56.180 ;
        RECT 137.290 -56.280 139.360 -56.270 ;
        RECT 140.830 -56.280 141.080 -56.190 ;
        RECT 141.940 -56.280 142.230 -56.230 ;
        RECT 137.290 -56.410 142.230 -56.280 ;
        RECT 137.290 -56.520 137.540 -56.410 ;
        RECT 139.040 -56.420 142.230 -56.410 ;
        RECT 139.040 -56.500 139.360 -56.420 ;
        RECT 140.830 -56.510 141.080 -56.420 ;
        RECT 141.940 -56.460 142.230 -56.420 ;
        RECT -39.900 -58.630 -39.580 -58.570 ;
        RECT -37.240 -58.620 -37.010 -58.590 ;
        RECT -33.190 -58.620 -32.960 -58.590 ;
        RECT -25.740 -58.620 -25.510 -58.590 ;
        RECT -21.690 -58.620 -21.460 -58.590 ;
        RECT -13.920 -58.620 -13.690 -58.590 ;
        RECT -9.870 -58.620 -9.640 -58.590 ;
        RECT -2.110 -58.620 -1.880 -58.590 ;
        RECT 1.940 -58.620 2.170 -58.590 ;
        RECT 9.700 -58.620 9.930 -58.590 ;
        RECT 13.750 -58.620 13.980 -58.590 ;
        RECT 21.520 -58.620 21.750 -58.590 ;
        RECT 25.570 -58.620 25.800 -58.590 ;
        RECT 33.340 -58.620 33.570 -58.590 ;
        RECT 37.390 -58.620 37.620 -58.590 ;
        RECT 45.160 -58.620 45.390 -58.590 ;
        RECT 49.210 -58.620 49.440 -58.590 ;
        RECT 56.980 -58.620 57.210 -58.590 ;
        RECT 61.030 -58.620 61.260 -58.590 ;
        RECT 68.800 -58.620 69.030 -58.590 ;
        RECT 72.850 -58.620 73.080 -58.590 ;
        RECT 80.620 -58.620 80.850 -58.590 ;
        RECT 84.670 -58.620 84.900 -58.590 ;
        RECT 92.460 -58.620 92.690 -58.590 ;
        RECT 96.510 -58.620 96.740 -58.590 ;
        RECT 104.300 -58.620 104.530 -58.590 ;
        RECT 108.350 -58.620 108.580 -58.590 ;
        RECT 116.170 -58.620 116.400 -58.590 ;
        RECT 120.220 -58.620 120.450 -58.590 ;
        RECT 128.040 -58.620 128.270 -58.590 ;
        RECT 132.090 -58.620 132.320 -58.590 ;
        RECT 137.050 -58.620 137.280 -58.590 ;
        RECT 141.100 -58.620 141.330 -58.590 ;
        RECT -37.290 -58.630 -36.960 -58.620 ;
        RECT -33.240 -58.630 -32.910 -58.620 ;
        RECT -25.790 -58.630 -25.460 -58.620 ;
        RECT -21.740 -58.630 -21.410 -58.620 ;
        RECT -13.970 -58.630 -13.640 -58.620 ;
        RECT -9.920 -58.630 -9.590 -58.620 ;
        RECT -2.160 -58.630 -1.830 -58.620 ;
        RECT 1.890 -58.630 2.220 -58.620 ;
        RECT 9.650 -58.630 9.980 -58.620 ;
        RECT 13.700 -58.630 14.030 -58.620 ;
        RECT 21.470 -58.630 21.800 -58.620 ;
        RECT 25.520 -58.630 25.850 -58.620 ;
        RECT 33.290 -58.630 33.620 -58.620 ;
        RECT 37.340 -58.630 37.670 -58.620 ;
        RECT 45.110 -58.630 45.440 -58.620 ;
        RECT 49.160 -58.630 49.490 -58.620 ;
        RECT 56.930 -58.630 57.260 -58.620 ;
        RECT 60.980 -58.630 61.310 -58.620 ;
        RECT 68.750 -58.630 69.080 -58.620 ;
        RECT 72.800 -58.630 73.130 -58.620 ;
        RECT 80.570 -58.630 80.900 -58.620 ;
        RECT 84.620 -58.630 84.950 -58.620 ;
        RECT 92.410 -58.630 92.740 -58.620 ;
        RECT 96.460 -58.630 96.790 -58.620 ;
        RECT 104.250 -58.630 104.580 -58.620 ;
        RECT 108.300 -58.630 108.630 -58.620 ;
        RECT 116.120 -58.630 116.450 -58.620 ;
        RECT 120.170 -58.630 120.500 -58.620 ;
        RECT 127.990 -58.630 128.320 -58.620 ;
        RECT 132.040 -58.630 132.370 -58.620 ;
        RECT 137.000 -58.630 137.330 -58.620 ;
        RECT 141.050 -58.630 141.380 -58.620 ;
        RECT -39.900 -58.780 142.470 -58.630 ;
        RECT -39.900 -58.830 -39.580 -58.780 ;
        RECT -37.290 -58.790 -36.960 -58.780 ;
        RECT -33.240 -58.790 -32.910 -58.780 ;
        RECT -25.790 -58.790 -25.460 -58.780 ;
        RECT -21.740 -58.790 -21.410 -58.780 ;
        RECT -13.970 -58.790 -13.640 -58.780 ;
        RECT -9.920 -58.790 -9.590 -58.780 ;
        RECT -2.160 -58.790 -1.830 -58.780 ;
        RECT 1.890 -58.790 2.220 -58.780 ;
        RECT 9.650 -58.790 9.980 -58.780 ;
        RECT 13.700 -58.790 14.030 -58.780 ;
        RECT 21.470 -58.790 21.800 -58.780 ;
        RECT 25.520 -58.790 25.850 -58.780 ;
        RECT 33.290 -58.790 33.620 -58.780 ;
        RECT 37.340 -58.790 37.670 -58.780 ;
        RECT 45.110 -58.790 45.440 -58.780 ;
        RECT 49.160 -58.790 49.490 -58.780 ;
        RECT 56.930 -58.790 57.260 -58.780 ;
        RECT 60.980 -58.790 61.310 -58.780 ;
        RECT 68.750 -58.790 69.080 -58.780 ;
        RECT 72.800 -58.790 73.130 -58.780 ;
        RECT 80.570 -58.790 80.900 -58.780 ;
        RECT 84.620 -58.790 84.950 -58.780 ;
        RECT 92.410 -58.790 92.740 -58.780 ;
        RECT 96.460 -58.790 96.790 -58.780 ;
        RECT 104.250 -58.790 104.580 -58.780 ;
        RECT 108.300 -58.790 108.630 -58.780 ;
        RECT 116.120 -58.790 116.450 -58.780 ;
        RECT 120.170 -58.790 120.500 -58.780 ;
        RECT 127.990 -58.790 128.320 -58.780 ;
        RECT 132.040 -58.790 132.370 -58.780 ;
        RECT 137.000 -58.790 137.330 -58.780 ;
        RECT 141.050 -58.790 141.380 -58.780 ;
        RECT -37.240 -58.820 -37.010 -58.790 ;
        RECT -33.190 -58.820 -32.960 -58.790 ;
        RECT -25.740 -58.820 -25.510 -58.790 ;
        RECT -21.690 -58.820 -21.460 -58.790 ;
        RECT -13.920 -58.820 -13.690 -58.790 ;
        RECT -9.870 -58.820 -9.640 -58.790 ;
        RECT -2.110 -58.820 -1.880 -58.790 ;
        RECT 1.940 -58.820 2.170 -58.790 ;
        RECT 9.700 -58.820 9.930 -58.790 ;
        RECT 13.750 -58.820 13.980 -58.790 ;
        RECT 21.520 -58.820 21.750 -58.790 ;
        RECT 25.570 -58.820 25.800 -58.790 ;
        RECT 33.340 -58.820 33.570 -58.790 ;
        RECT 37.390 -58.820 37.620 -58.790 ;
        RECT 45.160 -58.820 45.390 -58.790 ;
        RECT 49.210 -58.820 49.440 -58.790 ;
        RECT 56.980 -58.820 57.210 -58.790 ;
        RECT 61.030 -58.820 61.260 -58.790 ;
        RECT 68.800 -58.820 69.030 -58.790 ;
        RECT 72.850 -58.820 73.080 -58.790 ;
        RECT 80.620 -58.820 80.850 -58.790 ;
        RECT 84.670 -58.820 84.900 -58.790 ;
        RECT 92.460 -58.820 92.690 -58.790 ;
        RECT 96.510 -58.820 96.740 -58.790 ;
        RECT 104.300 -58.820 104.530 -58.790 ;
        RECT 108.350 -58.820 108.580 -58.790 ;
        RECT 116.170 -58.820 116.400 -58.790 ;
        RECT 120.220 -58.820 120.450 -58.790 ;
        RECT 128.040 -58.820 128.270 -58.790 ;
        RECT 132.090 -58.820 132.320 -58.790 ;
        RECT 137.050 -58.820 137.280 -58.790 ;
        RECT 141.100 -58.820 141.330 -58.790 ;
        RECT -37.000 -61.000 -36.750 -60.890 ;
        RECT -35.250 -60.990 -34.930 -60.910 ;
        RECT -33.460 -60.990 -33.210 -60.900 ;
        RECT -32.360 -60.990 -32.070 -60.940 ;
        RECT -35.250 -61.000 -32.070 -60.990 ;
        RECT -37.000 -61.130 -32.070 -61.000 ;
        RECT -37.000 -61.140 -34.930 -61.130 ;
        RECT -37.000 -61.250 -36.750 -61.140 ;
        RECT -35.250 -61.230 -34.930 -61.140 ;
        RECT -33.460 -61.220 -33.210 -61.130 ;
        RECT -32.360 -61.170 -32.070 -61.130 ;
        RECT -25.500 -61.000 -25.250 -60.890 ;
        RECT -23.750 -60.990 -23.430 -60.910 ;
        RECT -21.960 -60.990 -21.710 -60.900 ;
        RECT -20.860 -60.990 -20.570 -60.940 ;
        RECT -23.750 -61.000 -20.570 -60.990 ;
        RECT -25.500 -61.130 -20.570 -61.000 ;
        RECT -25.500 -61.140 -23.430 -61.130 ;
        RECT -25.500 -61.250 -25.250 -61.140 ;
        RECT -23.750 -61.230 -23.430 -61.140 ;
        RECT -21.960 -61.220 -21.710 -61.130 ;
        RECT -20.860 -61.170 -20.570 -61.130 ;
        RECT -13.680 -61.000 -13.430 -60.890 ;
        RECT -11.930 -60.990 -11.610 -60.910 ;
        RECT -10.140 -60.990 -9.890 -60.900 ;
        RECT -9.040 -60.990 -8.750 -60.940 ;
        RECT -11.930 -61.000 -8.750 -60.990 ;
        RECT -13.680 -61.130 -8.750 -61.000 ;
        RECT -13.680 -61.140 -11.610 -61.130 ;
        RECT -13.680 -61.250 -13.430 -61.140 ;
        RECT -11.930 -61.230 -11.610 -61.140 ;
        RECT -10.140 -61.220 -9.890 -61.130 ;
        RECT -9.040 -61.170 -8.750 -61.130 ;
        RECT -1.870 -61.000 -1.620 -60.890 ;
        RECT -0.120 -60.990 0.200 -60.910 ;
        RECT 1.670 -60.990 1.920 -60.900 ;
        RECT 2.770 -60.990 3.060 -60.940 ;
        RECT -0.120 -61.000 3.060 -60.990 ;
        RECT -1.870 -61.130 3.060 -61.000 ;
        RECT -1.870 -61.140 0.200 -61.130 ;
        RECT -1.870 -61.250 -1.620 -61.140 ;
        RECT -0.120 -61.230 0.200 -61.140 ;
        RECT 1.670 -61.220 1.920 -61.130 ;
        RECT 2.770 -61.170 3.060 -61.130 ;
        RECT 9.940 -61.000 10.190 -60.890 ;
        RECT 11.690 -60.990 12.010 -60.910 ;
        RECT 13.480 -60.990 13.730 -60.900 ;
        RECT 14.580 -60.990 14.870 -60.940 ;
        RECT 11.690 -61.000 14.870 -60.990 ;
        RECT 9.940 -61.130 14.870 -61.000 ;
        RECT 9.940 -61.140 12.010 -61.130 ;
        RECT 9.940 -61.250 10.190 -61.140 ;
        RECT 11.690 -61.230 12.010 -61.140 ;
        RECT 13.480 -61.220 13.730 -61.130 ;
        RECT 14.580 -61.170 14.870 -61.130 ;
        RECT 21.760 -61.000 22.010 -60.890 ;
        RECT 23.510 -60.990 23.830 -60.910 ;
        RECT 25.300 -60.990 25.550 -60.900 ;
        RECT 26.400 -60.990 26.690 -60.940 ;
        RECT 23.510 -61.000 26.690 -60.990 ;
        RECT 21.760 -61.130 26.690 -61.000 ;
        RECT 21.760 -61.140 23.830 -61.130 ;
        RECT 21.760 -61.250 22.010 -61.140 ;
        RECT 23.510 -61.230 23.830 -61.140 ;
        RECT 25.300 -61.220 25.550 -61.130 ;
        RECT 26.400 -61.170 26.690 -61.130 ;
        RECT 33.580 -61.000 33.830 -60.890 ;
        RECT 35.330 -60.990 35.650 -60.910 ;
        RECT 37.120 -60.990 37.370 -60.900 ;
        RECT 38.220 -60.990 38.510 -60.940 ;
        RECT 35.330 -61.000 38.510 -60.990 ;
        RECT 33.580 -61.130 38.510 -61.000 ;
        RECT 33.580 -61.140 35.650 -61.130 ;
        RECT 33.580 -61.250 33.830 -61.140 ;
        RECT 35.330 -61.230 35.650 -61.140 ;
        RECT 37.120 -61.220 37.370 -61.130 ;
        RECT 38.220 -61.170 38.510 -61.130 ;
        RECT 45.400 -61.000 45.650 -60.890 ;
        RECT 47.150 -60.990 47.470 -60.910 ;
        RECT 48.940 -60.990 49.190 -60.900 ;
        RECT 50.040 -60.990 50.330 -60.940 ;
        RECT 47.150 -61.000 50.330 -60.990 ;
        RECT 45.400 -61.130 50.330 -61.000 ;
        RECT 45.400 -61.140 47.470 -61.130 ;
        RECT 45.400 -61.250 45.650 -61.140 ;
        RECT 47.150 -61.230 47.470 -61.140 ;
        RECT 48.940 -61.220 49.190 -61.130 ;
        RECT 50.040 -61.170 50.330 -61.130 ;
        RECT 57.220 -61.000 57.470 -60.890 ;
        RECT 58.970 -60.990 59.290 -60.910 ;
        RECT 60.760 -60.990 61.010 -60.900 ;
        RECT 61.860 -60.990 62.150 -60.940 ;
        RECT 58.970 -61.000 62.150 -60.990 ;
        RECT 57.220 -61.130 62.150 -61.000 ;
        RECT 57.220 -61.140 59.290 -61.130 ;
        RECT 57.220 -61.250 57.470 -61.140 ;
        RECT 58.970 -61.230 59.290 -61.140 ;
        RECT 60.760 -61.220 61.010 -61.130 ;
        RECT 61.860 -61.170 62.150 -61.130 ;
        RECT 69.040 -61.000 69.290 -60.890 ;
        RECT 70.790 -60.990 71.110 -60.910 ;
        RECT 72.580 -60.990 72.830 -60.900 ;
        RECT 73.680 -60.990 73.970 -60.940 ;
        RECT 70.790 -61.000 73.970 -60.990 ;
        RECT 69.040 -61.130 73.970 -61.000 ;
        RECT 69.040 -61.140 71.110 -61.130 ;
        RECT 69.040 -61.250 69.290 -61.140 ;
        RECT 70.790 -61.230 71.110 -61.140 ;
        RECT 72.580 -61.220 72.830 -61.130 ;
        RECT 73.680 -61.170 73.970 -61.130 ;
        RECT 80.860 -61.000 81.110 -60.890 ;
        RECT 82.610 -60.990 82.930 -60.910 ;
        RECT 84.400 -60.990 84.650 -60.900 ;
        RECT 85.500 -60.990 85.790 -60.940 ;
        RECT 82.610 -61.000 85.790 -60.990 ;
        RECT 80.860 -61.130 85.790 -61.000 ;
        RECT 80.860 -61.140 82.930 -61.130 ;
        RECT 80.860 -61.250 81.110 -61.140 ;
        RECT 82.610 -61.230 82.930 -61.140 ;
        RECT 84.400 -61.220 84.650 -61.130 ;
        RECT 85.500 -61.170 85.790 -61.130 ;
        RECT 92.700 -61.000 92.950 -60.890 ;
        RECT 94.450 -60.990 94.770 -60.910 ;
        RECT 96.240 -60.990 96.490 -60.900 ;
        RECT 97.340 -60.990 97.630 -60.940 ;
        RECT 94.450 -61.000 97.630 -60.990 ;
        RECT 92.700 -61.130 97.630 -61.000 ;
        RECT 92.700 -61.140 94.770 -61.130 ;
        RECT 92.700 -61.250 92.950 -61.140 ;
        RECT 94.450 -61.230 94.770 -61.140 ;
        RECT 96.240 -61.220 96.490 -61.130 ;
        RECT 97.340 -61.170 97.630 -61.130 ;
        RECT 104.540 -61.000 104.790 -60.890 ;
        RECT 106.290 -60.990 106.610 -60.910 ;
        RECT 108.080 -60.990 108.330 -60.900 ;
        RECT 109.180 -60.990 109.470 -60.940 ;
        RECT 106.290 -61.000 109.470 -60.990 ;
        RECT 104.540 -61.130 109.470 -61.000 ;
        RECT 104.540 -61.140 106.610 -61.130 ;
        RECT 104.540 -61.250 104.790 -61.140 ;
        RECT 106.290 -61.230 106.610 -61.140 ;
        RECT 108.080 -61.220 108.330 -61.130 ;
        RECT 109.180 -61.170 109.470 -61.130 ;
        RECT 116.410 -61.000 116.660 -60.890 ;
        RECT 118.160 -60.990 118.480 -60.910 ;
        RECT 119.950 -60.990 120.200 -60.900 ;
        RECT 121.050 -60.990 121.340 -60.940 ;
        RECT 118.160 -61.000 121.340 -60.990 ;
        RECT 116.410 -61.130 121.340 -61.000 ;
        RECT 116.410 -61.140 118.480 -61.130 ;
        RECT 116.410 -61.250 116.660 -61.140 ;
        RECT 118.160 -61.230 118.480 -61.140 ;
        RECT 119.950 -61.220 120.200 -61.130 ;
        RECT 121.050 -61.170 121.340 -61.130 ;
        RECT 128.280 -61.000 128.530 -60.890 ;
        RECT 130.030 -60.990 130.350 -60.910 ;
        RECT 131.820 -60.990 132.070 -60.900 ;
        RECT 132.920 -60.990 133.210 -60.940 ;
        RECT 130.030 -61.000 133.210 -60.990 ;
        RECT 128.280 -61.130 133.210 -61.000 ;
        RECT 128.280 -61.140 130.350 -61.130 ;
        RECT 128.280 -61.250 128.530 -61.140 ;
        RECT 130.030 -61.230 130.350 -61.140 ;
        RECT 131.820 -61.220 132.070 -61.130 ;
        RECT 132.920 -61.170 133.210 -61.130 ;
        RECT 137.290 -61.000 137.540 -60.890 ;
        RECT 139.040 -60.990 139.360 -60.910 ;
        RECT 140.830 -60.990 141.080 -60.900 ;
        RECT 141.930 -60.990 142.220 -60.940 ;
        RECT 139.040 -61.000 142.220 -60.990 ;
        RECT 137.290 -61.130 142.220 -61.000 ;
        RECT 137.290 -61.140 139.360 -61.130 ;
        RECT 137.290 -61.250 137.540 -61.140 ;
        RECT 139.040 -61.230 139.360 -61.140 ;
        RECT 140.830 -61.220 141.080 -61.130 ;
        RECT 141.930 -61.170 142.220 -61.130 ;
        RECT -36.370 -63.230 -36.140 -63.160 ;
        RECT -30.700 -63.230 -30.380 -63.170 ;
        RECT -36.370 -63.370 -30.380 -63.230 ;
        RECT -36.370 -63.450 -36.140 -63.370 ;
        RECT -30.700 -63.430 -30.380 -63.370 ;
        RECT -24.930 -63.230 -24.630 -63.160 ;
        RECT -19.140 -63.230 -18.820 -63.170 ;
        RECT -24.930 -63.370 -18.820 -63.230 ;
        RECT -24.930 -63.450 -24.630 -63.370 ;
        RECT -19.140 -63.430 -18.820 -63.370 ;
        RECT -13.110 -63.230 -12.820 -63.160 ;
        RECT -7.450 -63.230 -7.130 -63.170 ;
        RECT -13.110 -63.370 -7.130 -63.230 ;
        RECT -13.110 -63.450 -12.820 -63.370 ;
        RECT -7.450 -63.430 -7.130 -63.370 ;
        RECT -1.360 -63.230 -1.070 -63.160 ;
        RECT 4.460 -63.230 4.780 -63.170 ;
        RECT -1.360 -63.370 4.780 -63.230 ;
        RECT -1.360 -63.440 -1.070 -63.370 ;
        RECT 4.460 -63.430 4.780 -63.370 ;
        RECT 10.520 -63.230 10.810 -63.160 ;
        RECT 16.230 -63.230 16.550 -63.170 ;
        RECT 10.520 -63.370 16.550 -63.230 ;
        RECT 10.520 -63.450 10.810 -63.370 ;
        RECT 16.230 -63.430 16.550 -63.370 ;
        RECT 22.360 -63.230 22.650 -63.160 ;
        RECT 28.000 -63.230 28.320 -63.170 ;
        RECT 22.360 -63.370 28.320 -63.230 ;
        RECT 22.360 -63.450 22.650 -63.370 ;
        RECT 28.000 -63.430 28.320 -63.370 ;
        RECT 34.070 -63.230 34.360 -63.160 ;
        RECT 39.820 -63.230 40.140 -63.170 ;
        RECT 34.070 -63.370 40.140 -63.230 ;
        RECT 34.070 -63.450 34.360 -63.370 ;
        RECT 39.820 -63.430 40.140 -63.370 ;
        RECT 45.940 -63.230 46.230 -63.160 ;
        RECT 51.680 -63.230 52.000 -63.170 ;
        RECT 45.940 -63.370 52.000 -63.230 ;
        RECT 45.940 -63.450 46.230 -63.370 ;
        RECT 51.680 -63.430 52.000 -63.370 ;
        RECT 57.820 -63.230 58.110 -63.160 ;
        RECT 63.470 -63.230 63.790 -63.170 ;
        RECT 57.820 -63.370 63.790 -63.230 ;
        RECT 57.820 -63.450 58.110 -63.370 ;
        RECT 63.470 -63.430 63.790 -63.370 ;
        RECT 69.490 -63.230 69.780 -63.160 ;
        RECT 75.350 -63.230 75.670 -63.170 ;
        RECT 69.490 -63.370 75.670 -63.230 ;
        RECT 69.490 -63.450 69.780 -63.370 ;
        RECT 75.350 -63.430 75.670 -63.370 ;
        RECT 81.310 -63.230 81.600 -63.160 ;
        RECT 87.080 -63.230 87.400 -63.170 ;
        RECT 81.310 -63.370 87.400 -63.230 ;
        RECT 81.310 -63.450 81.600 -63.370 ;
        RECT 87.080 -63.430 87.400 -63.370 ;
        RECT 93.170 -63.230 93.460 -63.160 ;
        RECT 98.900 -63.230 99.220 -63.170 ;
        RECT 93.170 -63.370 99.220 -63.230 ;
        RECT 93.170 -63.450 93.460 -63.370 ;
        RECT 98.900 -63.430 99.220 -63.370 ;
        RECT 104.930 -63.230 105.220 -63.160 ;
        RECT 110.790 -63.230 111.110 -63.170 ;
        RECT 104.930 -63.370 111.110 -63.230 ;
        RECT 104.930 -63.450 105.220 -63.370 ;
        RECT 110.790 -63.430 111.110 -63.370 ;
        RECT 116.720 -63.230 117.010 -63.160 ;
        RECT 122.740 -63.230 123.060 -63.170 ;
        RECT 116.720 -63.370 123.060 -63.230 ;
        RECT 116.720 -63.450 117.010 -63.370 ;
        RECT 122.740 -63.430 123.060 -63.370 ;
        RECT 128.740 -63.230 129.030 -63.160 ;
        RECT 134.500 -63.230 134.820 -63.170 ;
        RECT 128.740 -63.370 134.820 -63.230 ;
        RECT 128.740 -63.450 129.030 -63.370 ;
        RECT 134.500 -63.430 134.820 -63.370 ;
        RECT 137.730 -63.230 138.020 -63.160 ;
        RECT 143.540 -63.230 143.860 -63.170 ;
        RECT 137.730 -63.370 143.860 -63.230 ;
        RECT 137.730 -63.450 138.020 -63.370 ;
        RECT 143.540 -63.430 143.860 -63.370 ;
        RECT -40.570 -63.670 -40.250 -63.610 ;
        RECT -36.790 -63.670 -36.460 -63.620 ;
        RECT -33.720 -63.670 -33.390 -63.610 ;
        RECT -25.290 -63.670 -24.960 -63.620 ;
        RECT -22.220 -63.670 -21.890 -63.610 ;
        RECT -13.470 -63.670 -13.140 -63.620 ;
        RECT -10.400 -63.670 -10.070 -63.610 ;
        RECT -1.660 -63.670 -1.330 -63.620 ;
        RECT 1.410 -63.670 1.740 -63.610 ;
        RECT 10.150 -63.670 10.480 -63.620 ;
        RECT 13.220 -63.670 13.550 -63.610 ;
        RECT 21.970 -63.670 22.300 -63.620 ;
        RECT 25.040 -63.670 25.370 -63.610 ;
        RECT 33.790 -63.670 34.120 -63.620 ;
        RECT 36.860 -63.670 37.190 -63.610 ;
        RECT 45.610 -63.670 45.940 -63.620 ;
        RECT 48.680 -63.670 49.010 -63.610 ;
        RECT 57.430 -63.670 57.760 -63.620 ;
        RECT 60.500 -63.670 60.830 -63.610 ;
        RECT 69.250 -63.670 69.580 -63.620 ;
        RECT 72.320 -63.670 72.650 -63.610 ;
        RECT 81.070 -63.670 81.400 -63.620 ;
        RECT 84.140 -63.670 84.470 -63.610 ;
        RECT 92.910 -63.670 93.240 -63.620 ;
        RECT 95.980 -63.670 96.310 -63.610 ;
        RECT 104.750 -63.670 105.080 -63.620 ;
        RECT 107.820 -63.670 108.150 -63.610 ;
        RECT 116.620 -63.670 116.950 -63.620 ;
        RECT 119.690 -63.670 120.020 -63.610 ;
        RECT 128.490 -63.670 128.820 -63.620 ;
        RECT 131.560 -63.670 131.890 -63.610 ;
        RECT 137.500 -63.670 137.830 -63.620 ;
        RECT 140.570 -63.670 140.900 -63.610 ;
        RECT -40.570 -63.810 50.580 -63.670 ;
        RECT 50.850 -63.810 142.470 -63.670 ;
        RECT -40.570 -63.870 -40.250 -63.810 ;
        RECT -36.790 -63.860 -36.460 -63.810 ;
        RECT -33.720 -63.850 -33.390 -63.810 ;
        RECT -25.290 -63.860 -24.960 -63.810 ;
        RECT -22.220 -63.850 -21.890 -63.810 ;
        RECT -13.470 -63.860 -13.140 -63.810 ;
        RECT -10.400 -63.850 -10.070 -63.810 ;
        RECT -1.660 -63.860 -1.330 -63.810 ;
        RECT 1.410 -63.850 1.740 -63.810 ;
        RECT 10.150 -63.860 10.480 -63.810 ;
        RECT 13.220 -63.850 13.550 -63.810 ;
        RECT 21.970 -63.860 22.300 -63.810 ;
        RECT 25.040 -63.850 25.370 -63.810 ;
        RECT 33.790 -63.860 34.120 -63.810 ;
        RECT 36.860 -63.850 37.190 -63.810 ;
        RECT 45.610 -63.860 45.940 -63.810 ;
        RECT 48.680 -63.850 49.010 -63.810 ;
        RECT 57.430 -63.860 57.760 -63.810 ;
        RECT 60.500 -63.850 60.830 -63.810 ;
        RECT 69.250 -63.860 69.580 -63.810 ;
        RECT 72.320 -63.850 72.650 -63.810 ;
        RECT 81.070 -63.860 81.400 -63.810 ;
        RECT 84.140 -63.850 84.470 -63.810 ;
        RECT 92.910 -63.860 93.240 -63.810 ;
        RECT 95.980 -63.850 96.310 -63.810 ;
        RECT 104.750 -63.860 105.080 -63.810 ;
        RECT 107.820 -63.850 108.150 -63.810 ;
        RECT 116.620 -63.860 116.950 -63.810 ;
        RECT 119.690 -63.850 120.020 -63.810 ;
        RECT 128.490 -63.860 128.820 -63.810 ;
        RECT 131.560 -63.850 131.890 -63.810 ;
        RECT 137.500 -63.860 137.830 -63.810 ;
        RECT 140.570 -63.850 140.900 -63.810 ;
        RECT -41.230 -64.070 -40.910 -64.010 ;
        RECT -37.860 -64.040 -37.570 -64.010 ;
        RECT -37.900 -64.070 -37.570 -64.040 ;
        RECT -32.640 -64.060 -32.350 -64.030 ;
        RECT -26.360 -64.040 -26.070 -64.010 ;
        RECT -32.640 -64.070 -32.310 -64.060 ;
        RECT -26.400 -64.070 -26.070 -64.040 ;
        RECT -21.140 -64.060 -20.850 -64.030 ;
        RECT -14.540 -64.040 -14.250 -64.010 ;
        RECT -21.140 -64.070 -20.810 -64.060 ;
        RECT -14.580 -64.070 -14.250 -64.040 ;
        RECT -9.320 -64.060 -9.030 -64.030 ;
        RECT -2.730 -64.040 -2.440 -64.010 ;
        RECT -9.320 -64.070 -8.990 -64.060 ;
        RECT -2.770 -64.070 -2.440 -64.040 ;
        RECT 2.490 -64.060 2.780 -64.030 ;
        RECT 9.080 -64.040 9.370 -64.010 ;
        RECT 2.490 -64.070 2.820 -64.060 ;
        RECT 9.040 -64.070 9.370 -64.040 ;
        RECT 14.300 -64.060 14.590 -64.030 ;
        RECT 20.900 -64.040 21.190 -64.010 ;
        RECT 14.300 -64.070 14.630 -64.060 ;
        RECT 20.860 -64.070 21.190 -64.040 ;
        RECT 26.120 -64.060 26.410 -64.030 ;
        RECT 32.720 -64.040 33.010 -64.010 ;
        RECT 26.120 -64.070 26.450 -64.060 ;
        RECT 32.680 -64.070 33.010 -64.040 ;
        RECT 37.940 -64.060 38.230 -64.030 ;
        RECT 44.540 -64.040 44.830 -64.010 ;
        RECT 37.940 -64.070 38.270 -64.060 ;
        RECT 44.500 -64.070 44.830 -64.040 ;
        RECT 49.760 -64.060 50.050 -64.030 ;
        RECT 56.360 -64.040 56.650 -64.010 ;
        RECT 49.760 -64.070 50.090 -64.060 ;
        RECT 56.320 -64.070 56.650 -64.040 ;
        RECT 61.580 -64.060 61.870 -64.030 ;
        RECT 68.180 -64.040 68.470 -64.010 ;
        RECT 61.580 -64.070 61.910 -64.060 ;
        RECT 68.140 -64.070 68.470 -64.040 ;
        RECT 73.400 -64.060 73.690 -64.030 ;
        RECT 80.000 -64.040 80.290 -64.010 ;
        RECT 73.400 -64.070 73.730 -64.060 ;
        RECT 79.960 -64.070 80.290 -64.040 ;
        RECT 85.220 -64.060 85.510 -64.030 ;
        RECT 91.840 -64.040 92.130 -64.010 ;
        RECT 85.220 -64.070 85.550 -64.060 ;
        RECT 91.800 -64.070 92.130 -64.040 ;
        RECT 97.060 -64.060 97.350 -64.030 ;
        RECT 103.680 -64.040 103.970 -64.010 ;
        RECT 97.060 -64.070 97.390 -64.060 ;
        RECT 103.640 -64.070 103.970 -64.040 ;
        RECT 108.900 -64.060 109.190 -64.030 ;
        RECT 115.550 -64.040 115.840 -64.010 ;
        RECT 108.900 -64.070 109.230 -64.060 ;
        RECT 115.510 -64.070 115.840 -64.040 ;
        RECT 120.770 -64.060 121.060 -64.030 ;
        RECT 127.420 -64.040 127.710 -64.010 ;
        RECT 120.770 -64.070 121.100 -64.060 ;
        RECT 127.380 -64.070 127.710 -64.040 ;
        RECT 132.640 -64.060 132.930 -64.030 ;
        RECT 136.430 -64.040 136.720 -64.010 ;
        RECT 132.640 -64.070 132.970 -64.060 ;
        RECT 136.390 -64.070 136.720 -64.040 ;
        RECT 141.650 -64.060 141.940 -64.030 ;
        RECT 141.650 -64.070 141.980 -64.060 ;
        RECT -41.230 -64.210 50.580 -64.070 ;
        RECT 50.850 -64.210 142.470 -64.070 ;
        RECT -41.230 -64.270 -40.910 -64.210 ;
        RECT -37.900 -64.220 -37.570 -64.210 ;
        RECT -37.860 -64.250 -37.570 -64.220 ;
        RECT -32.640 -64.240 -32.310 -64.210 ;
        RECT -26.400 -64.220 -26.070 -64.210 ;
        RECT -32.640 -64.270 -32.350 -64.240 ;
        RECT -26.360 -64.250 -26.070 -64.220 ;
        RECT -21.140 -64.240 -20.810 -64.210 ;
        RECT -14.580 -64.220 -14.250 -64.210 ;
        RECT -21.140 -64.270 -20.850 -64.240 ;
        RECT -14.540 -64.250 -14.250 -64.220 ;
        RECT -9.320 -64.240 -8.990 -64.210 ;
        RECT -2.770 -64.220 -2.440 -64.210 ;
        RECT -9.320 -64.270 -9.030 -64.240 ;
        RECT -2.730 -64.250 -2.440 -64.220 ;
        RECT 2.490 -64.240 2.820 -64.210 ;
        RECT 9.040 -64.220 9.370 -64.210 ;
        RECT 2.490 -64.270 2.780 -64.240 ;
        RECT 9.080 -64.250 9.370 -64.220 ;
        RECT 14.300 -64.240 14.630 -64.210 ;
        RECT 20.860 -64.220 21.190 -64.210 ;
        RECT 14.300 -64.270 14.590 -64.240 ;
        RECT 20.900 -64.250 21.190 -64.220 ;
        RECT 26.120 -64.240 26.450 -64.210 ;
        RECT 32.680 -64.220 33.010 -64.210 ;
        RECT 26.120 -64.270 26.410 -64.240 ;
        RECT 32.720 -64.250 33.010 -64.220 ;
        RECT 37.940 -64.240 38.270 -64.210 ;
        RECT 44.500 -64.220 44.830 -64.210 ;
        RECT 37.940 -64.270 38.230 -64.240 ;
        RECT 44.540 -64.250 44.830 -64.220 ;
        RECT 49.760 -64.240 50.090 -64.210 ;
        RECT 56.320 -64.220 56.650 -64.210 ;
        RECT 49.760 -64.270 50.050 -64.240 ;
        RECT 56.360 -64.250 56.650 -64.220 ;
        RECT 61.580 -64.240 61.910 -64.210 ;
        RECT 68.140 -64.220 68.470 -64.210 ;
        RECT 61.580 -64.270 61.870 -64.240 ;
        RECT 68.180 -64.250 68.470 -64.220 ;
        RECT 73.400 -64.240 73.730 -64.210 ;
        RECT 79.960 -64.220 80.290 -64.210 ;
        RECT 73.400 -64.270 73.690 -64.240 ;
        RECT 80.000 -64.250 80.290 -64.220 ;
        RECT 85.220 -64.240 85.550 -64.210 ;
        RECT 91.800 -64.220 92.130 -64.210 ;
        RECT 85.220 -64.270 85.510 -64.240 ;
        RECT 91.840 -64.250 92.130 -64.220 ;
        RECT 97.060 -64.240 97.390 -64.210 ;
        RECT 103.640 -64.220 103.970 -64.210 ;
        RECT 97.060 -64.270 97.350 -64.240 ;
        RECT 103.680 -64.250 103.970 -64.220 ;
        RECT 108.900 -64.240 109.230 -64.210 ;
        RECT 115.510 -64.220 115.840 -64.210 ;
        RECT 108.900 -64.270 109.190 -64.240 ;
        RECT 115.550 -64.250 115.840 -64.220 ;
        RECT 120.770 -64.240 121.100 -64.210 ;
        RECT 127.380 -64.220 127.710 -64.210 ;
        RECT 120.770 -64.270 121.060 -64.240 ;
        RECT 127.420 -64.250 127.710 -64.220 ;
        RECT 132.640 -64.240 132.970 -64.210 ;
        RECT 136.390 -64.220 136.720 -64.210 ;
        RECT 132.640 -64.270 132.930 -64.240 ;
        RECT 136.430 -64.250 136.720 -64.220 ;
        RECT 141.650 -64.240 141.980 -64.210 ;
        RECT 141.650 -64.270 141.940 -64.240 ;
        RECT -37.940 -64.700 -37.650 -64.640 ;
        RECT -36.460 -64.700 -36.170 -64.610 ;
        RECT -37.940 -64.840 -36.170 -64.700 ;
        RECT -37.940 -64.890 -37.650 -64.840 ;
        RECT -36.460 -64.860 -36.170 -64.840 ;
        RECT -34.010 -64.670 -33.720 -64.600 ;
        RECT -32.560 -64.670 -32.270 -64.630 ;
        RECT -34.010 -64.810 -32.270 -64.670 ;
        RECT -34.010 -64.850 -33.720 -64.810 ;
        RECT -32.560 -64.880 -32.270 -64.810 ;
        RECT -26.440 -64.700 -26.150 -64.640 ;
        RECT -24.960 -64.700 -24.670 -64.610 ;
        RECT -26.440 -64.840 -24.670 -64.700 ;
        RECT -26.440 -64.890 -26.150 -64.840 ;
        RECT -24.960 -64.860 -24.670 -64.840 ;
        RECT -22.510 -64.670 -22.220 -64.600 ;
        RECT -21.060 -64.670 -20.770 -64.630 ;
        RECT -22.510 -64.810 -20.770 -64.670 ;
        RECT -22.510 -64.850 -22.220 -64.810 ;
        RECT -21.060 -64.880 -20.770 -64.810 ;
        RECT -14.620 -64.700 -14.330 -64.640 ;
        RECT -13.140 -64.700 -12.850 -64.610 ;
        RECT -14.620 -64.840 -12.850 -64.700 ;
        RECT -14.620 -64.890 -14.330 -64.840 ;
        RECT -13.140 -64.860 -12.850 -64.840 ;
        RECT -10.690 -64.670 -10.400 -64.600 ;
        RECT -9.240 -64.670 -8.950 -64.630 ;
        RECT -10.690 -64.810 -8.950 -64.670 ;
        RECT -10.690 -64.850 -10.400 -64.810 ;
        RECT -9.240 -64.880 -8.950 -64.810 ;
        RECT -2.810 -64.700 -2.520 -64.640 ;
        RECT -1.330 -64.700 -1.040 -64.610 ;
        RECT -2.810 -64.840 -1.040 -64.700 ;
        RECT -2.810 -64.890 -2.520 -64.840 ;
        RECT -1.330 -64.860 -1.040 -64.840 ;
        RECT 1.120 -64.670 1.410 -64.600 ;
        RECT 2.570 -64.670 2.860 -64.630 ;
        RECT 1.120 -64.810 2.860 -64.670 ;
        RECT 1.120 -64.850 1.410 -64.810 ;
        RECT 2.570 -64.880 2.860 -64.810 ;
        RECT 9.000 -64.700 9.290 -64.640 ;
        RECT 10.480 -64.700 10.770 -64.610 ;
        RECT 9.000 -64.840 10.770 -64.700 ;
        RECT 9.000 -64.890 9.290 -64.840 ;
        RECT 10.480 -64.860 10.770 -64.840 ;
        RECT 12.930 -64.670 13.220 -64.600 ;
        RECT 14.380 -64.670 14.670 -64.630 ;
        RECT 12.930 -64.810 14.670 -64.670 ;
        RECT 12.930 -64.850 13.220 -64.810 ;
        RECT 14.380 -64.880 14.670 -64.810 ;
        RECT 20.820 -64.700 21.110 -64.640 ;
        RECT 22.300 -64.700 22.590 -64.610 ;
        RECT 20.820 -64.840 22.590 -64.700 ;
        RECT 20.820 -64.890 21.110 -64.840 ;
        RECT 22.300 -64.860 22.590 -64.840 ;
        RECT 24.750 -64.670 25.040 -64.600 ;
        RECT 26.200 -64.670 26.490 -64.630 ;
        RECT 24.750 -64.810 26.490 -64.670 ;
        RECT 24.750 -64.850 25.040 -64.810 ;
        RECT 26.200 -64.880 26.490 -64.810 ;
        RECT 32.640 -64.700 32.930 -64.640 ;
        RECT 34.120 -64.700 34.410 -64.610 ;
        RECT 32.640 -64.840 34.410 -64.700 ;
        RECT 32.640 -64.890 32.930 -64.840 ;
        RECT 34.120 -64.860 34.410 -64.840 ;
        RECT 36.570 -64.670 36.860 -64.600 ;
        RECT 38.020 -64.670 38.310 -64.630 ;
        RECT 36.570 -64.810 38.310 -64.670 ;
        RECT 36.570 -64.850 36.860 -64.810 ;
        RECT 38.020 -64.880 38.310 -64.810 ;
        RECT 44.460 -64.700 44.750 -64.640 ;
        RECT 45.940 -64.700 46.230 -64.610 ;
        RECT 44.460 -64.840 46.230 -64.700 ;
        RECT 44.460 -64.890 44.750 -64.840 ;
        RECT 45.940 -64.860 46.230 -64.840 ;
        RECT 48.390 -64.670 48.680 -64.600 ;
        RECT 49.840 -64.670 50.130 -64.630 ;
        RECT 48.390 -64.810 50.130 -64.670 ;
        RECT 48.390 -64.850 48.680 -64.810 ;
        RECT 49.840 -64.880 50.130 -64.810 ;
        RECT 56.280 -64.700 56.570 -64.640 ;
        RECT 57.760 -64.700 58.050 -64.610 ;
        RECT 56.280 -64.840 58.050 -64.700 ;
        RECT 56.280 -64.890 56.570 -64.840 ;
        RECT 57.760 -64.860 58.050 -64.840 ;
        RECT 60.210 -64.670 60.500 -64.600 ;
        RECT 61.660 -64.670 61.950 -64.630 ;
        RECT 60.210 -64.810 61.950 -64.670 ;
        RECT 60.210 -64.850 60.500 -64.810 ;
        RECT 61.660 -64.880 61.950 -64.810 ;
        RECT 68.100 -64.700 68.390 -64.640 ;
        RECT 69.580 -64.700 69.870 -64.610 ;
        RECT 68.100 -64.840 69.870 -64.700 ;
        RECT 68.100 -64.890 68.390 -64.840 ;
        RECT 69.580 -64.860 69.870 -64.840 ;
        RECT 72.030 -64.670 72.320 -64.600 ;
        RECT 73.480 -64.670 73.770 -64.630 ;
        RECT 72.030 -64.810 73.770 -64.670 ;
        RECT 72.030 -64.850 72.320 -64.810 ;
        RECT 73.480 -64.880 73.770 -64.810 ;
        RECT 79.920 -64.700 80.210 -64.640 ;
        RECT 81.400 -64.700 81.690 -64.610 ;
        RECT 79.920 -64.840 81.690 -64.700 ;
        RECT 79.920 -64.890 80.210 -64.840 ;
        RECT 81.400 -64.860 81.690 -64.840 ;
        RECT 83.850 -64.670 84.140 -64.600 ;
        RECT 85.300 -64.670 85.590 -64.630 ;
        RECT 83.850 -64.810 85.590 -64.670 ;
        RECT 83.850 -64.850 84.140 -64.810 ;
        RECT 85.300 -64.880 85.590 -64.810 ;
        RECT 91.760 -64.700 92.050 -64.640 ;
        RECT 93.240 -64.700 93.530 -64.610 ;
        RECT 91.760 -64.840 93.530 -64.700 ;
        RECT 91.760 -64.890 92.050 -64.840 ;
        RECT 93.240 -64.860 93.530 -64.840 ;
        RECT 95.690 -64.670 95.980 -64.600 ;
        RECT 97.140 -64.670 97.430 -64.630 ;
        RECT 95.690 -64.810 97.430 -64.670 ;
        RECT 95.690 -64.850 95.980 -64.810 ;
        RECT 97.140 -64.880 97.430 -64.810 ;
        RECT 103.600 -64.700 103.890 -64.640 ;
        RECT 105.080 -64.700 105.370 -64.610 ;
        RECT 103.600 -64.840 105.370 -64.700 ;
        RECT 103.600 -64.890 103.890 -64.840 ;
        RECT 105.080 -64.860 105.370 -64.840 ;
        RECT 107.530 -64.670 107.820 -64.600 ;
        RECT 108.980 -64.670 109.270 -64.630 ;
        RECT 107.530 -64.810 109.270 -64.670 ;
        RECT 107.530 -64.850 107.820 -64.810 ;
        RECT 108.980 -64.880 109.270 -64.810 ;
        RECT 115.470 -64.700 115.760 -64.640 ;
        RECT 116.950 -64.700 117.240 -64.610 ;
        RECT 115.470 -64.840 117.240 -64.700 ;
        RECT 115.470 -64.890 115.760 -64.840 ;
        RECT 116.950 -64.860 117.240 -64.840 ;
        RECT 119.400 -64.670 119.690 -64.600 ;
        RECT 120.850 -64.670 121.140 -64.630 ;
        RECT 119.400 -64.810 121.140 -64.670 ;
        RECT 119.400 -64.850 119.690 -64.810 ;
        RECT 120.850 -64.880 121.140 -64.810 ;
        RECT 127.340 -64.700 127.630 -64.640 ;
        RECT 128.820 -64.700 129.110 -64.610 ;
        RECT 127.340 -64.840 129.110 -64.700 ;
        RECT 127.340 -64.890 127.630 -64.840 ;
        RECT 128.820 -64.860 129.110 -64.840 ;
        RECT 131.270 -64.670 131.560 -64.600 ;
        RECT 132.720 -64.670 133.010 -64.630 ;
        RECT 131.270 -64.810 133.010 -64.670 ;
        RECT 131.270 -64.850 131.560 -64.810 ;
        RECT 132.720 -64.880 133.010 -64.810 ;
        RECT 136.350 -64.700 136.640 -64.640 ;
        RECT 137.830 -64.700 138.120 -64.610 ;
        RECT 136.350 -64.840 138.120 -64.700 ;
        RECT 136.350 -64.890 136.640 -64.840 ;
        RECT 137.830 -64.860 138.120 -64.840 ;
        RECT 140.280 -64.670 140.570 -64.600 ;
        RECT 141.730 -64.670 142.020 -64.630 ;
        RECT 140.280 -64.810 142.020 -64.670 ;
        RECT 140.280 -64.850 140.570 -64.810 ;
        RECT 141.730 -64.880 142.020 -64.810 ;
        RECT -36.460 -65.370 -36.170 -65.320 ;
        RECT -35.500 -65.370 -35.210 -65.320 ;
        RECT -36.460 -65.510 -35.210 -65.370 ;
        RECT -36.460 -65.570 -36.170 -65.510 ;
        RECT -35.500 -65.570 -35.210 -65.510 ;
        RECT -24.960 -65.370 -24.670 -65.320 ;
        RECT -24.000 -65.370 -23.710 -65.320 ;
        RECT -24.960 -65.510 -23.710 -65.370 ;
        RECT -24.960 -65.570 -24.670 -65.510 ;
        RECT -24.000 -65.570 -23.710 -65.510 ;
        RECT -13.140 -65.370 -12.850 -65.320 ;
        RECT -12.180 -65.370 -11.890 -65.320 ;
        RECT -13.140 -65.510 -11.890 -65.370 ;
        RECT -13.140 -65.570 -12.850 -65.510 ;
        RECT -12.180 -65.570 -11.890 -65.510 ;
        RECT -1.330 -65.370 -1.040 -65.320 ;
        RECT -0.370 -65.370 -0.080 -65.320 ;
        RECT -1.330 -65.510 -0.080 -65.370 ;
        RECT -1.330 -65.570 -1.040 -65.510 ;
        RECT -0.370 -65.570 -0.080 -65.510 ;
        RECT 10.480 -65.370 10.770 -65.320 ;
        RECT 11.440 -65.370 11.730 -65.320 ;
        RECT 10.480 -65.510 11.730 -65.370 ;
        RECT 10.480 -65.570 10.770 -65.510 ;
        RECT 11.440 -65.570 11.730 -65.510 ;
        RECT 22.300 -65.370 22.590 -65.320 ;
        RECT 23.260 -65.370 23.550 -65.320 ;
        RECT 22.300 -65.510 23.550 -65.370 ;
        RECT 22.300 -65.570 22.590 -65.510 ;
        RECT 23.260 -65.570 23.550 -65.510 ;
        RECT 34.120 -65.370 34.410 -65.320 ;
        RECT 35.080 -65.370 35.370 -65.320 ;
        RECT 34.120 -65.510 35.370 -65.370 ;
        RECT 34.120 -65.570 34.410 -65.510 ;
        RECT 35.080 -65.570 35.370 -65.510 ;
        RECT 45.940 -65.370 46.230 -65.320 ;
        RECT 46.900 -65.370 47.190 -65.320 ;
        RECT 45.940 -65.510 47.190 -65.370 ;
        RECT 45.940 -65.570 46.230 -65.510 ;
        RECT 46.900 -65.570 47.190 -65.510 ;
        RECT 57.760 -65.370 58.050 -65.320 ;
        RECT 58.720 -65.370 59.010 -65.320 ;
        RECT 57.760 -65.510 59.010 -65.370 ;
        RECT 57.760 -65.570 58.050 -65.510 ;
        RECT 58.720 -65.570 59.010 -65.510 ;
        RECT 69.580 -65.370 69.870 -65.320 ;
        RECT 70.540 -65.370 70.830 -65.320 ;
        RECT 69.580 -65.510 70.830 -65.370 ;
        RECT 69.580 -65.570 69.870 -65.510 ;
        RECT 70.540 -65.570 70.830 -65.510 ;
        RECT 81.400 -65.370 81.690 -65.320 ;
        RECT 82.360 -65.370 82.650 -65.320 ;
        RECT 81.400 -65.510 82.650 -65.370 ;
        RECT 81.400 -65.570 81.690 -65.510 ;
        RECT 82.360 -65.570 82.650 -65.510 ;
        RECT 93.240 -65.370 93.530 -65.320 ;
        RECT 94.200 -65.370 94.490 -65.320 ;
        RECT 93.240 -65.510 94.490 -65.370 ;
        RECT 93.240 -65.570 93.530 -65.510 ;
        RECT 94.200 -65.570 94.490 -65.510 ;
        RECT 105.080 -65.370 105.370 -65.320 ;
        RECT 106.040 -65.370 106.330 -65.320 ;
        RECT 105.080 -65.510 106.330 -65.370 ;
        RECT 105.080 -65.570 105.370 -65.510 ;
        RECT 106.040 -65.570 106.330 -65.510 ;
        RECT 116.950 -65.370 117.240 -65.320 ;
        RECT 117.910 -65.370 118.200 -65.320 ;
        RECT 116.950 -65.510 118.200 -65.370 ;
        RECT 116.950 -65.570 117.240 -65.510 ;
        RECT 117.910 -65.570 118.200 -65.510 ;
        RECT 128.820 -65.370 129.110 -65.320 ;
        RECT 129.780 -65.370 130.070 -65.320 ;
        RECT 128.820 -65.510 130.070 -65.370 ;
        RECT 128.820 -65.570 129.110 -65.510 ;
        RECT 129.780 -65.570 130.070 -65.510 ;
        RECT 137.830 -65.370 138.120 -65.320 ;
        RECT 138.790 -65.370 139.080 -65.320 ;
        RECT 137.830 -65.510 139.080 -65.370 ;
        RECT 137.830 -65.570 138.120 -65.510 ;
        RECT 138.790 -65.570 139.080 -65.510 ;
        RECT -37.860 -66.040 -37.620 -66.030 ;
        RECT -26.360 -66.040 -26.120 -66.030 ;
        RECT -14.540 -66.040 -14.300 -66.030 ;
        RECT -2.730 -66.040 -2.490 -66.030 ;
        RECT 9.080 -66.040 9.320 -66.030 ;
        RECT 20.900 -66.040 21.140 -66.030 ;
        RECT 32.720 -66.040 32.960 -66.030 ;
        RECT 44.540 -66.040 44.780 -66.030 ;
        RECT 56.360 -66.040 56.600 -66.030 ;
        RECT 68.180 -66.040 68.420 -66.030 ;
        RECT 80.000 -66.040 80.240 -66.030 ;
        RECT 91.840 -66.040 92.080 -66.030 ;
        RECT 103.680 -66.040 103.920 -66.030 ;
        RECT 115.550 -66.040 115.790 -66.030 ;
        RECT 127.420 -66.040 127.660 -66.030 ;
        RECT 136.430 -66.040 136.670 -66.030 ;
        RECT -37.900 -66.360 -37.580 -66.040 ;
        RECT -34.970 -66.180 -34.680 -66.130 ;
        RECT -34.010 -66.180 -33.720 -66.140 ;
        RECT -34.970 -66.320 -33.720 -66.180 ;
        RECT -34.970 -66.380 -34.680 -66.320 ;
        RECT -34.010 -66.390 -33.720 -66.320 ;
        RECT -26.400 -66.360 -26.080 -66.040 ;
        RECT -23.470 -66.180 -23.180 -66.130 ;
        RECT -22.510 -66.180 -22.220 -66.140 ;
        RECT -23.470 -66.320 -22.220 -66.180 ;
        RECT -23.470 -66.380 -23.180 -66.320 ;
        RECT -22.510 -66.390 -22.220 -66.320 ;
        RECT -14.580 -66.360 -14.260 -66.040 ;
        RECT -11.650 -66.180 -11.360 -66.130 ;
        RECT -10.690 -66.180 -10.400 -66.140 ;
        RECT -11.650 -66.320 -10.400 -66.180 ;
        RECT -11.650 -66.380 -11.360 -66.320 ;
        RECT -10.690 -66.390 -10.400 -66.320 ;
        RECT -2.770 -66.360 -2.450 -66.040 ;
        RECT 0.160 -66.180 0.450 -66.130 ;
        RECT 1.120 -66.180 1.410 -66.140 ;
        RECT 0.160 -66.320 1.410 -66.180 ;
        RECT 0.160 -66.380 0.450 -66.320 ;
        RECT 1.120 -66.390 1.410 -66.320 ;
        RECT 9.040 -66.360 9.360 -66.040 ;
        RECT 11.970 -66.180 12.260 -66.130 ;
        RECT 12.930 -66.180 13.220 -66.140 ;
        RECT 11.970 -66.320 13.220 -66.180 ;
        RECT 11.970 -66.380 12.260 -66.320 ;
        RECT 12.930 -66.390 13.220 -66.320 ;
        RECT 20.860 -66.360 21.180 -66.040 ;
        RECT 23.790 -66.180 24.080 -66.130 ;
        RECT 24.750 -66.180 25.040 -66.140 ;
        RECT 23.790 -66.320 25.040 -66.180 ;
        RECT 23.790 -66.380 24.080 -66.320 ;
        RECT 24.750 -66.390 25.040 -66.320 ;
        RECT 32.680 -66.360 33.000 -66.040 ;
        RECT 35.610 -66.180 35.900 -66.130 ;
        RECT 36.570 -66.180 36.860 -66.140 ;
        RECT 35.610 -66.320 36.860 -66.180 ;
        RECT 35.610 -66.380 35.900 -66.320 ;
        RECT 36.570 -66.390 36.860 -66.320 ;
        RECT 44.500 -66.360 44.820 -66.040 ;
        RECT 47.430 -66.180 47.720 -66.130 ;
        RECT 48.390 -66.180 48.680 -66.140 ;
        RECT 47.430 -66.320 48.680 -66.180 ;
        RECT 47.430 -66.380 47.720 -66.320 ;
        RECT 48.390 -66.390 48.680 -66.320 ;
        RECT 56.320 -66.360 56.640 -66.040 ;
        RECT 59.250 -66.180 59.540 -66.130 ;
        RECT 60.210 -66.180 60.500 -66.140 ;
        RECT 59.250 -66.320 60.500 -66.180 ;
        RECT 59.250 -66.380 59.540 -66.320 ;
        RECT 60.210 -66.390 60.500 -66.320 ;
        RECT 68.140 -66.360 68.460 -66.040 ;
        RECT 71.070 -66.180 71.360 -66.130 ;
        RECT 72.030 -66.180 72.320 -66.140 ;
        RECT 71.070 -66.320 72.320 -66.180 ;
        RECT 71.070 -66.380 71.360 -66.320 ;
        RECT 72.030 -66.390 72.320 -66.320 ;
        RECT 79.960 -66.360 80.280 -66.040 ;
        RECT 82.890 -66.180 83.180 -66.130 ;
        RECT 83.850 -66.180 84.140 -66.140 ;
        RECT 82.890 -66.320 84.140 -66.180 ;
        RECT 82.890 -66.380 83.180 -66.320 ;
        RECT 83.850 -66.390 84.140 -66.320 ;
        RECT 91.800 -66.360 92.120 -66.040 ;
        RECT 94.730 -66.180 95.020 -66.130 ;
        RECT 95.690 -66.180 95.980 -66.140 ;
        RECT 94.730 -66.320 95.980 -66.180 ;
        RECT 94.730 -66.380 95.020 -66.320 ;
        RECT 95.690 -66.390 95.980 -66.320 ;
        RECT 103.640 -66.360 103.960 -66.040 ;
        RECT 106.570 -66.180 106.860 -66.130 ;
        RECT 107.530 -66.180 107.820 -66.140 ;
        RECT 106.570 -66.320 107.820 -66.180 ;
        RECT 106.570 -66.380 106.860 -66.320 ;
        RECT 107.530 -66.390 107.820 -66.320 ;
        RECT 115.510 -66.360 115.830 -66.040 ;
        RECT 118.440 -66.180 118.730 -66.130 ;
        RECT 119.400 -66.180 119.690 -66.140 ;
        RECT 118.440 -66.320 119.690 -66.180 ;
        RECT 118.440 -66.380 118.730 -66.320 ;
        RECT 119.400 -66.390 119.690 -66.320 ;
        RECT 127.380 -66.360 127.700 -66.040 ;
        RECT 130.310 -66.180 130.600 -66.130 ;
        RECT 131.270 -66.180 131.560 -66.140 ;
        RECT 130.310 -66.320 131.560 -66.180 ;
        RECT 130.310 -66.380 130.600 -66.320 ;
        RECT 131.270 -66.390 131.560 -66.320 ;
        RECT 136.390 -66.360 136.710 -66.040 ;
        RECT 139.320 -66.180 139.610 -66.130 ;
        RECT 140.280 -66.180 140.570 -66.140 ;
        RECT 139.320 -66.320 140.570 -66.180 ;
        RECT 139.320 -66.380 139.610 -66.320 ;
        RECT 140.280 -66.390 140.570 -66.320 ;
        RECT -38.290 -66.920 -38.000 -66.870 ;
        RECT -36.900 -66.920 -36.610 -66.870 ;
        RECT -38.290 -67.060 -36.610 -66.920 ;
        RECT -38.290 -67.120 -38.000 -67.060 ;
        RECT -36.900 -67.120 -36.610 -67.060 ;
        RECT -33.570 -66.920 -33.280 -66.860 ;
        RECT -32.210 -66.920 -31.920 -66.870 ;
        RECT -33.570 -67.060 -31.920 -66.920 ;
        RECT -33.570 -67.110 -33.280 -67.060 ;
        RECT -32.210 -67.120 -31.920 -67.060 ;
        RECT -26.790 -66.920 -26.500 -66.870 ;
        RECT -25.400 -66.920 -25.110 -66.870 ;
        RECT -26.790 -67.060 -25.110 -66.920 ;
        RECT -26.790 -67.120 -26.500 -67.060 ;
        RECT -25.400 -67.120 -25.110 -67.060 ;
        RECT -22.070 -66.920 -21.780 -66.860 ;
        RECT -20.710 -66.920 -20.420 -66.870 ;
        RECT -22.070 -67.060 -20.420 -66.920 ;
        RECT -22.070 -67.110 -21.780 -67.060 ;
        RECT -20.710 -67.120 -20.420 -67.060 ;
        RECT -14.970 -66.920 -14.680 -66.870 ;
        RECT -13.580 -66.920 -13.290 -66.870 ;
        RECT -14.970 -67.060 -13.290 -66.920 ;
        RECT -14.970 -67.120 -14.680 -67.060 ;
        RECT -13.580 -67.120 -13.290 -67.060 ;
        RECT -10.250 -66.920 -9.960 -66.860 ;
        RECT -8.890 -66.920 -8.600 -66.870 ;
        RECT -10.250 -67.060 -8.600 -66.920 ;
        RECT -10.250 -67.110 -9.960 -67.060 ;
        RECT -8.890 -67.120 -8.600 -67.060 ;
        RECT -3.160 -66.920 -2.870 -66.870 ;
        RECT -1.770 -66.920 -1.480 -66.870 ;
        RECT -3.160 -67.060 -1.480 -66.920 ;
        RECT -3.160 -67.120 -2.870 -67.060 ;
        RECT -1.770 -67.120 -1.480 -67.060 ;
        RECT 1.560 -66.920 1.850 -66.860 ;
        RECT 2.920 -66.920 3.210 -66.870 ;
        RECT 1.560 -67.060 3.210 -66.920 ;
        RECT 1.560 -67.110 1.850 -67.060 ;
        RECT 2.920 -67.120 3.210 -67.060 ;
        RECT 8.650 -66.920 8.940 -66.870 ;
        RECT 10.040 -66.920 10.330 -66.870 ;
        RECT 8.650 -67.060 10.330 -66.920 ;
        RECT 8.650 -67.120 8.940 -67.060 ;
        RECT 10.040 -67.120 10.330 -67.060 ;
        RECT 13.370 -66.920 13.660 -66.860 ;
        RECT 14.730 -66.920 15.020 -66.870 ;
        RECT 13.370 -67.060 15.020 -66.920 ;
        RECT 13.370 -67.110 13.660 -67.060 ;
        RECT 14.730 -67.120 15.020 -67.060 ;
        RECT 20.470 -66.920 20.760 -66.870 ;
        RECT 21.860 -66.920 22.150 -66.870 ;
        RECT 20.470 -67.060 22.150 -66.920 ;
        RECT 20.470 -67.120 20.760 -67.060 ;
        RECT 21.860 -67.120 22.150 -67.060 ;
        RECT 25.190 -66.920 25.480 -66.860 ;
        RECT 26.550 -66.920 26.840 -66.870 ;
        RECT 25.190 -67.060 26.840 -66.920 ;
        RECT 25.190 -67.110 25.480 -67.060 ;
        RECT 26.550 -67.120 26.840 -67.060 ;
        RECT 32.290 -66.920 32.580 -66.870 ;
        RECT 33.680 -66.920 33.970 -66.870 ;
        RECT 32.290 -67.060 33.970 -66.920 ;
        RECT 32.290 -67.120 32.580 -67.060 ;
        RECT 33.680 -67.120 33.970 -67.060 ;
        RECT 37.010 -66.920 37.300 -66.860 ;
        RECT 38.370 -66.920 38.660 -66.870 ;
        RECT 37.010 -67.060 38.660 -66.920 ;
        RECT 37.010 -67.110 37.300 -67.060 ;
        RECT 38.370 -67.120 38.660 -67.060 ;
        RECT 44.110 -66.920 44.400 -66.870 ;
        RECT 45.500 -66.920 45.790 -66.870 ;
        RECT 44.110 -67.060 45.790 -66.920 ;
        RECT 44.110 -67.120 44.400 -67.060 ;
        RECT 45.500 -67.120 45.790 -67.060 ;
        RECT 48.830 -66.920 49.120 -66.860 ;
        RECT 50.190 -66.920 50.480 -66.870 ;
        RECT 48.830 -67.060 50.480 -66.920 ;
        RECT 48.830 -67.110 49.120 -67.060 ;
        RECT 50.190 -67.120 50.480 -67.060 ;
        RECT 55.930 -66.920 56.220 -66.870 ;
        RECT 57.320 -66.920 57.610 -66.870 ;
        RECT 55.930 -67.060 57.610 -66.920 ;
        RECT 55.930 -67.120 56.220 -67.060 ;
        RECT 57.320 -67.120 57.610 -67.060 ;
        RECT 60.650 -66.920 60.940 -66.860 ;
        RECT 62.010 -66.920 62.300 -66.870 ;
        RECT 60.650 -67.060 62.300 -66.920 ;
        RECT 60.650 -67.110 60.940 -67.060 ;
        RECT 62.010 -67.120 62.300 -67.060 ;
        RECT 67.750 -66.920 68.040 -66.870 ;
        RECT 69.140 -66.920 69.430 -66.870 ;
        RECT 67.750 -67.060 69.430 -66.920 ;
        RECT 67.750 -67.120 68.040 -67.060 ;
        RECT 69.140 -67.120 69.430 -67.060 ;
        RECT 72.470 -66.920 72.760 -66.860 ;
        RECT 73.830 -66.920 74.120 -66.870 ;
        RECT 72.470 -67.060 74.120 -66.920 ;
        RECT 72.470 -67.110 72.760 -67.060 ;
        RECT 73.830 -67.120 74.120 -67.060 ;
        RECT 79.570 -66.920 79.860 -66.870 ;
        RECT 80.960 -66.920 81.250 -66.870 ;
        RECT 79.570 -67.060 81.250 -66.920 ;
        RECT 79.570 -67.120 79.860 -67.060 ;
        RECT 80.960 -67.120 81.250 -67.060 ;
        RECT 84.290 -66.920 84.580 -66.860 ;
        RECT 85.650 -66.920 85.940 -66.870 ;
        RECT 84.290 -67.060 85.940 -66.920 ;
        RECT 84.290 -67.110 84.580 -67.060 ;
        RECT 85.650 -67.120 85.940 -67.060 ;
        RECT 91.410 -66.920 91.700 -66.870 ;
        RECT 92.800 -66.920 93.090 -66.870 ;
        RECT 91.410 -67.060 93.090 -66.920 ;
        RECT 91.410 -67.120 91.700 -67.060 ;
        RECT 92.800 -67.120 93.090 -67.060 ;
        RECT 96.130 -66.920 96.420 -66.860 ;
        RECT 97.490 -66.920 97.780 -66.870 ;
        RECT 96.130 -67.060 97.780 -66.920 ;
        RECT 96.130 -67.110 96.420 -67.060 ;
        RECT 97.490 -67.120 97.780 -67.060 ;
        RECT 103.250 -66.920 103.540 -66.870 ;
        RECT 104.640 -66.920 104.930 -66.870 ;
        RECT 103.250 -67.060 104.930 -66.920 ;
        RECT 103.250 -67.120 103.540 -67.060 ;
        RECT 104.640 -67.120 104.930 -67.060 ;
        RECT 107.970 -66.920 108.260 -66.860 ;
        RECT 109.330 -66.920 109.620 -66.870 ;
        RECT 107.970 -67.060 109.620 -66.920 ;
        RECT 107.970 -67.110 108.260 -67.060 ;
        RECT 109.330 -67.120 109.620 -67.060 ;
        RECT 115.120 -66.920 115.410 -66.870 ;
        RECT 116.510 -66.920 116.800 -66.870 ;
        RECT 115.120 -67.060 116.800 -66.920 ;
        RECT 115.120 -67.120 115.410 -67.060 ;
        RECT 116.510 -67.120 116.800 -67.060 ;
        RECT 119.840 -66.920 120.130 -66.860 ;
        RECT 121.200 -66.920 121.490 -66.870 ;
        RECT 119.840 -67.060 121.490 -66.920 ;
        RECT 119.840 -67.110 120.130 -67.060 ;
        RECT 121.200 -67.120 121.490 -67.060 ;
        RECT 126.990 -66.920 127.280 -66.870 ;
        RECT 128.380 -66.920 128.670 -66.870 ;
        RECT 126.990 -67.060 128.670 -66.920 ;
        RECT 126.990 -67.120 127.280 -67.060 ;
        RECT 128.380 -67.120 128.670 -67.060 ;
        RECT 131.710 -66.920 132.000 -66.860 ;
        RECT 133.070 -66.920 133.360 -66.870 ;
        RECT 131.710 -67.060 133.360 -66.920 ;
        RECT 131.710 -67.110 132.000 -67.060 ;
        RECT 133.070 -67.120 133.360 -67.060 ;
        RECT 136.000 -66.920 136.290 -66.870 ;
        RECT 137.390 -66.920 137.680 -66.870 ;
        RECT 136.000 -67.060 137.680 -66.920 ;
        RECT 136.000 -67.120 136.290 -67.060 ;
        RECT 137.390 -67.120 137.680 -67.060 ;
        RECT 140.720 -66.920 141.010 -66.860 ;
        RECT 142.080 -66.920 142.370 -66.870 ;
        RECT 140.720 -67.060 142.370 -66.920 ;
        RECT 140.720 -67.110 141.010 -67.060 ;
        RECT 142.080 -67.120 142.370 -67.060 ;
        RECT -37.870 -68.630 -37.630 -68.620 ;
        RECT -26.370 -68.630 -26.130 -68.620 ;
        RECT -14.550 -68.630 -14.310 -68.620 ;
        RECT -2.740 -68.630 -2.500 -68.620 ;
        RECT 9.070 -68.630 9.310 -68.620 ;
        RECT 20.890 -68.630 21.130 -68.620 ;
        RECT 32.710 -68.630 32.950 -68.620 ;
        RECT 44.530 -68.630 44.770 -68.620 ;
        RECT 56.350 -68.630 56.590 -68.620 ;
        RECT 68.170 -68.630 68.410 -68.620 ;
        RECT 79.990 -68.630 80.230 -68.620 ;
        RECT 91.830 -68.630 92.070 -68.620 ;
        RECT 103.670 -68.630 103.910 -68.620 ;
        RECT 115.540 -68.630 115.780 -68.620 ;
        RECT 127.410 -68.630 127.650 -68.620 ;
        RECT 136.420 -68.630 136.660 -68.620 ;
        RECT -37.910 -68.950 -37.590 -68.630 ;
        RECT -26.410 -68.950 -26.090 -68.630 ;
        RECT -14.590 -68.950 -14.270 -68.630 ;
        RECT -2.780 -68.950 -2.460 -68.630 ;
        RECT 9.030 -68.950 9.350 -68.630 ;
        RECT 20.850 -68.950 21.170 -68.630 ;
        RECT 32.670 -68.950 32.990 -68.630 ;
        RECT 44.490 -68.950 44.810 -68.630 ;
        RECT 56.310 -68.950 56.630 -68.630 ;
        RECT 68.130 -68.950 68.450 -68.630 ;
        RECT 79.950 -68.950 80.270 -68.630 ;
        RECT 91.790 -68.950 92.110 -68.630 ;
        RECT 103.630 -68.950 103.950 -68.630 ;
        RECT 115.500 -68.950 115.820 -68.630 ;
        RECT 127.370 -68.950 127.690 -68.630 ;
        RECT 136.380 -68.950 136.700 -68.630 ;
        RECT -39.160 -70.850 -38.840 -70.790 ;
        RECT -37.490 -70.850 -37.210 -70.780 ;
        RECT -33.000 -70.850 -32.680 -70.790 ;
        RECT -25.990 -70.850 -25.710 -70.780 ;
        RECT -21.500 -70.850 -21.180 -70.790 ;
        RECT -14.170 -70.850 -13.890 -70.780 ;
        RECT -9.680 -70.850 -9.360 -70.790 ;
        RECT -2.360 -70.850 -2.080 -70.780 ;
        RECT 2.130 -70.850 2.450 -70.790 ;
        RECT 9.450 -70.850 9.730 -70.780 ;
        RECT 13.940 -70.850 14.260 -70.790 ;
        RECT 21.270 -70.850 21.550 -70.780 ;
        RECT 25.760 -70.850 26.080 -70.790 ;
        RECT 33.090 -70.850 33.370 -70.780 ;
        RECT 37.580 -70.850 37.900 -70.790 ;
        RECT 44.910 -70.850 45.190 -70.780 ;
        RECT 49.400 -70.850 49.720 -70.790 ;
        RECT 56.730 -70.850 57.010 -70.780 ;
        RECT 61.220 -70.850 61.540 -70.790 ;
        RECT 68.550 -70.850 68.830 -70.780 ;
        RECT 73.040 -70.850 73.360 -70.790 ;
        RECT 80.370 -70.850 80.650 -70.780 ;
        RECT 84.860 -70.850 85.180 -70.790 ;
        RECT 92.210 -70.850 92.490 -70.780 ;
        RECT 96.700 -70.850 97.020 -70.790 ;
        RECT 104.050 -70.850 104.330 -70.780 ;
        RECT 108.540 -70.850 108.860 -70.790 ;
        RECT 115.920 -70.850 116.200 -70.780 ;
        RECT 120.410 -70.850 120.730 -70.790 ;
        RECT 127.790 -70.850 128.070 -70.780 ;
        RECT 132.280 -70.850 132.600 -70.790 ;
        RECT 136.800 -70.850 137.080 -70.780 ;
        RECT 141.290 -70.850 141.610 -70.790 ;
        RECT -39.160 -70.990 142.470 -70.850 ;
        RECT -39.160 -71.050 -38.840 -70.990 ;
        RECT -37.490 -71.080 -37.210 -70.990 ;
        RECT -33.000 -71.050 -32.680 -70.990 ;
        RECT -25.990 -71.080 -25.710 -70.990 ;
        RECT -21.500 -71.050 -21.180 -70.990 ;
        RECT -14.170 -71.080 -13.890 -70.990 ;
        RECT -9.680 -71.050 -9.360 -70.990 ;
        RECT -2.360 -71.080 -2.080 -70.990 ;
        RECT 2.130 -71.050 2.450 -70.990 ;
        RECT 9.450 -71.080 9.730 -70.990 ;
        RECT 13.940 -71.050 14.260 -70.990 ;
        RECT 21.270 -71.080 21.550 -70.990 ;
        RECT 25.760 -71.050 26.080 -70.990 ;
        RECT 33.090 -71.080 33.370 -70.990 ;
        RECT 37.580 -71.050 37.900 -70.990 ;
        RECT 44.910 -71.080 45.190 -70.990 ;
        RECT 49.400 -71.050 49.720 -70.990 ;
        RECT 56.730 -71.080 57.010 -70.990 ;
        RECT 61.220 -71.050 61.540 -70.990 ;
        RECT 68.550 -71.080 68.830 -70.990 ;
        RECT 73.040 -71.050 73.360 -70.990 ;
        RECT 80.370 -71.080 80.650 -70.990 ;
        RECT 84.860 -71.050 85.180 -70.990 ;
        RECT 92.210 -71.080 92.490 -70.990 ;
        RECT 96.700 -71.050 97.020 -70.990 ;
        RECT 104.050 -71.080 104.330 -70.990 ;
        RECT 108.540 -71.050 108.860 -70.990 ;
        RECT 115.920 -71.080 116.200 -70.990 ;
        RECT 120.410 -71.050 120.730 -70.990 ;
        RECT 127.790 -71.080 128.070 -70.990 ;
        RECT 132.280 -71.050 132.600 -70.990 ;
        RECT 136.800 -71.080 137.080 -70.990 ;
        RECT 141.290 -71.050 141.610 -70.990 ;
        RECT -32.210 -71.760 -31.920 -71.740 ;
        RECT -20.710 -71.760 -20.420 -71.730 ;
        RECT -8.890 -71.760 -8.600 -71.730 ;
        RECT 2.920 -71.760 3.210 -71.730 ;
        RECT 14.730 -71.760 15.020 -71.730 ;
        RECT 26.550 -71.760 26.840 -71.730 ;
        RECT 38.370 -71.760 38.660 -71.730 ;
        RECT 50.190 -71.760 50.480 -71.730 ;
        RECT 62.010 -71.760 62.300 -71.730 ;
        RECT 73.830 -71.760 74.120 -71.730 ;
        RECT 85.650 -71.760 85.940 -71.730 ;
        RECT 97.490 -71.760 97.780 -71.730 ;
        RECT 109.330 -71.760 109.620 -71.730 ;
        RECT 121.200 -71.760 121.490 -71.730 ;
        RECT 133.070 -71.760 133.360 -71.730 ;
        RECT 142.080 -71.760 142.370 -71.730 ;
        RECT 145.530 -71.760 145.850 -71.710 ;
        RECT -32.210 -71.930 145.850 -71.760 ;
        RECT -32.210 -71.970 -31.920 -71.930 ;
        RECT -20.710 -71.960 -20.420 -71.930 ;
        RECT -8.890 -71.960 -8.600 -71.930 ;
        RECT 2.920 -71.960 3.210 -71.930 ;
        RECT 14.730 -71.960 15.020 -71.930 ;
        RECT 26.550 -71.960 26.840 -71.930 ;
        RECT 38.370 -71.960 38.660 -71.930 ;
        RECT 50.190 -71.960 50.480 -71.930 ;
        RECT 62.010 -71.960 62.300 -71.930 ;
        RECT 73.830 -71.960 74.120 -71.930 ;
        RECT 85.650 -71.960 85.940 -71.930 ;
        RECT 97.490 -71.960 97.780 -71.930 ;
        RECT 109.330 -71.960 109.620 -71.930 ;
        RECT 121.200 -71.960 121.490 -71.930 ;
        RECT 133.070 -71.960 133.360 -71.930 ;
        RECT 142.080 -71.960 142.370 -71.930 ;
        RECT 145.530 -71.970 145.850 -71.930 ;
        RECT -32.990 -72.300 -32.640 -72.220 ;
        RECT -21.490 -72.300 -21.140 -72.220 ;
        RECT -9.670 -72.300 -9.320 -72.220 ;
        RECT 2.140 -72.300 2.490 -72.220 ;
        RECT 13.950 -72.300 14.300 -72.220 ;
        RECT 25.770 -72.300 26.120 -72.220 ;
        RECT 37.590 -72.300 37.940 -72.220 ;
        RECT 49.410 -72.300 49.760 -72.220 ;
        RECT 61.230 -72.300 61.580 -72.220 ;
        RECT 73.050 -72.300 73.400 -72.220 ;
        RECT 84.870 -72.300 85.220 -72.220 ;
        RECT 96.710 -72.300 97.060 -72.220 ;
        RECT 108.550 -72.300 108.900 -72.220 ;
        RECT 120.420 -72.300 120.770 -72.220 ;
        RECT 132.290 -72.300 132.640 -72.220 ;
        RECT 141.300 -72.300 141.650 -72.220 ;
        RECT -32.990 -72.560 -32.620 -72.300 ;
        RECT -21.490 -72.560 -21.120 -72.300 ;
        RECT -9.670 -72.560 -9.300 -72.300 ;
        RECT 2.140 -72.560 2.510 -72.300 ;
        RECT 13.950 -72.560 14.320 -72.300 ;
        RECT 25.770 -72.560 26.140 -72.300 ;
        RECT 37.590 -72.560 37.960 -72.300 ;
        RECT 49.410 -72.560 49.780 -72.300 ;
        RECT 61.230 -72.560 61.600 -72.300 ;
        RECT 73.050 -72.560 73.420 -72.300 ;
        RECT 84.870 -72.560 85.240 -72.300 ;
        RECT 96.710 -72.560 97.080 -72.300 ;
        RECT 108.550 -72.560 108.920 -72.300 ;
        RECT 120.420 -72.560 120.790 -72.300 ;
        RECT 132.290 -72.560 132.660 -72.300 ;
        RECT 141.300 -72.560 141.670 -72.300 ;
        RECT -32.210 -72.730 -31.920 -72.710 ;
        RECT -20.710 -72.730 -20.420 -72.700 ;
        RECT -8.890 -72.730 -8.600 -72.700 ;
        RECT 2.920 -72.730 3.210 -72.700 ;
        RECT 14.730 -72.730 15.020 -72.700 ;
        RECT 26.550 -72.730 26.840 -72.700 ;
        RECT 38.370 -72.730 38.660 -72.700 ;
        RECT 50.190 -72.730 50.480 -72.700 ;
        RECT 62.010 -72.730 62.300 -72.700 ;
        RECT 73.830 -72.730 74.120 -72.700 ;
        RECT 85.650 -72.730 85.940 -72.700 ;
        RECT 97.490 -72.730 97.780 -72.700 ;
        RECT 109.330 -72.730 109.620 -72.700 ;
        RECT 121.200 -72.730 121.490 -72.700 ;
        RECT 133.070 -72.730 133.360 -72.700 ;
        RECT 142.110 -72.730 142.340 -72.670 ;
        RECT 146.080 -72.730 146.400 -72.680 ;
        RECT -32.210 -72.900 146.400 -72.730 ;
        RECT -32.210 -72.940 -31.920 -72.900 ;
        RECT -20.710 -72.930 -20.420 -72.900 ;
        RECT -8.890 -72.930 -8.600 -72.900 ;
        RECT 2.920 -72.930 3.210 -72.900 ;
        RECT 14.730 -72.930 15.020 -72.900 ;
        RECT 26.550 -72.930 26.840 -72.900 ;
        RECT 38.370 -72.930 38.660 -72.900 ;
        RECT 50.190 -72.930 50.480 -72.900 ;
        RECT 62.010 -72.930 62.300 -72.900 ;
        RECT 73.830 -72.930 74.120 -72.900 ;
        RECT 85.650 -72.930 85.940 -72.900 ;
        RECT 97.490 -72.930 97.780 -72.900 ;
        RECT 109.330 -72.930 109.620 -72.900 ;
        RECT 121.200 -72.930 121.490 -72.900 ;
        RECT 133.070 -72.930 133.360 -72.900 ;
        RECT 142.110 -72.960 142.340 -72.900 ;
        RECT 146.080 -72.940 146.400 -72.900 ;
        RECT -39.130 -73.750 -38.870 -73.660 ;
        RECT -37.490 -73.750 -37.210 -73.660 ;
        RECT -33.000 -73.750 -32.680 -73.660 ;
        RECT -25.990 -73.750 -25.710 -73.660 ;
        RECT -21.500 -73.750 -21.180 -73.660 ;
        RECT -14.170 -73.750 -13.890 -73.660 ;
        RECT -9.680 -73.750 -9.360 -73.660 ;
        RECT -2.360 -73.750 -2.080 -73.660 ;
        RECT 2.130 -73.750 2.450 -73.660 ;
        RECT 9.450 -73.750 9.730 -73.660 ;
        RECT 13.940 -73.750 14.260 -73.660 ;
        RECT 21.270 -73.750 21.550 -73.660 ;
        RECT 25.760 -73.750 26.080 -73.660 ;
        RECT 33.090 -73.750 33.370 -73.660 ;
        RECT 37.580 -73.750 37.900 -73.660 ;
        RECT 44.910 -73.750 45.190 -73.660 ;
        RECT 49.400 -73.750 49.720 -73.660 ;
        RECT 56.730 -73.750 57.010 -73.660 ;
        RECT 61.220 -73.750 61.540 -73.660 ;
        RECT 68.550 -73.750 68.830 -73.660 ;
        RECT 73.040 -73.750 73.360 -73.660 ;
        RECT 80.370 -73.750 80.650 -73.660 ;
        RECT 84.860 -73.750 85.180 -73.660 ;
        RECT 92.210 -73.750 92.490 -73.660 ;
        RECT 96.700 -73.750 97.020 -73.660 ;
        RECT 104.050 -73.750 104.330 -73.660 ;
        RECT 108.540 -73.750 108.860 -73.660 ;
        RECT 115.920 -73.750 116.200 -73.660 ;
        RECT 120.410 -73.750 120.730 -73.660 ;
        RECT 127.790 -73.750 128.070 -73.660 ;
        RECT 132.280 -73.750 132.600 -73.660 ;
        RECT 136.800 -73.750 137.080 -73.660 ;
        RECT 141.290 -73.750 141.610 -73.660 ;
        RECT -39.130 -73.890 142.470 -73.750 ;
        RECT -39.130 -73.980 -38.870 -73.890 ;
        RECT -37.490 -73.960 -37.210 -73.890 ;
        RECT -33.000 -73.980 -32.680 -73.890 ;
        RECT -25.990 -73.960 -25.710 -73.890 ;
        RECT -21.500 -73.980 -21.180 -73.890 ;
        RECT -14.170 -73.960 -13.890 -73.890 ;
        RECT -9.680 -73.980 -9.360 -73.890 ;
        RECT -2.360 -73.960 -2.080 -73.890 ;
        RECT 2.130 -73.980 2.450 -73.890 ;
        RECT 9.450 -73.960 9.730 -73.890 ;
        RECT 13.940 -73.980 14.260 -73.890 ;
        RECT 21.270 -73.960 21.550 -73.890 ;
        RECT 25.760 -73.980 26.080 -73.890 ;
        RECT 33.090 -73.960 33.370 -73.890 ;
        RECT 37.580 -73.980 37.900 -73.890 ;
        RECT 44.910 -73.960 45.190 -73.890 ;
        RECT 49.400 -73.980 49.720 -73.890 ;
        RECT 56.730 -73.960 57.010 -73.890 ;
        RECT 61.220 -73.980 61.540 -73.890 ;
        RECT 68.550 -73.960 68.830 -73.890 ;
        RECT 73.040 -73.980 73.360 -73.890 ;
        RECT 80.370 -73.960 80.650 -73.890 ;
        RECT 84.860 -73.980 85.180 -73.890 ;
        RECT 92.210 -73.960 92.490 -73.890 ;
        RECT 96.700 -73.980 97.020 -73.890 ;
        RECT 104.050 -73.960 104.330 -73.890 ;
        RECT 108.540 -73.980 108.860 -73.890 ;
        RECT 115.920 -73.960 116.200 -73.890 ;
        RECT 120.410 -73.980 120.730 -73.890 ;
        RECT 127.790 -73.960 128.070 -73.890 ;
        RECT 132.280 -73.980 132.600 -73.890 ;
        RECT 136.800 -73.960 137.080 -73.890 ;
        RECT 141.290 -73.980 141.610 -73.890 ;
        RECT -37.870 -75.800 -37.630 -75.790 ;
        RECT -26.370 -75.800 -26.130 -75.790 ;
        RECT -14.550 -75.800 -14.310 -75.790 ;
        RECT -2.740 -75.800 -2.500 -75.790 ;
        RECT 9.070 -75.800 9.310 -75.790 ;
        RECT 20.890 -75.800 21.130 -75.790 ;
        RECT 32.710 -75.800 32.950 -75.790 ;
        RECT 44.530 -75.800 44.770 -75.790 ;
        RECT 56.350 -75.800 56.590 -75.790 ;
        RECT 68.170 -75.800 68.410 -75.790 ;
        RECT 79.990 -75.800 80.230 -75.790 ;
        RECT 91.830 -75.800 92.070 -75.790 ;
        RECT 103.670 -75.800 103.910 -75.790 ;
        RECT 115.540 -75.800 115.780 -75.790 ;
        RECT 127.410 -75.800 127.650 -75.790 ;
        RECT 136.420 -75.800 136.660 -75.790 ;
        RECT -37.910 -76.120 -37.590 -75.800 ;
        RECT -26.410 -76.120 -26.090 -75.800 ;
        RECT -14.590 -76.120 -14.270 -75.800 ;
        RECT -2.780 -76.120 -2.460 -75.800 ;
        RECT 9.030 -76.120 9.350 -75.800 ;
        RECT 20.850 -76.120 21.170 -75.800 ;
        RECT 32.670 -76.120 32.990 -75.800 ;
        RECT 44.490 -76.120 44.810 -75.800 ;
        RECT 56.310 -76.120 56.630 -75.800 ;
        RECT 68.130 -76.120 68.450 -75.800 ;
        RECT 79.950 -76.120 80.270 -75.800 ;
        RECT 91.790 -76.120 92.110 -75.800 ;
        RECT 103.630 -76.120 103.950 -75.800 ;
        RECT 115.500 -76.120 115.820 -75.800 ;
        RECT 127.370 -76.120 127.690 -75.800 ;
        RECT 136.380 -76.120 136.700 -75.800 ;
        RECT -38.290 -77.680 -38.000 -77.620 ;
        RECT -36.900 -77.680 -36.610 -77.620 ;
        RECT -38.290 -77.820 -36.610 -77.680 ;
        RECT -38.290 -77.870 -38.000 -77.820 ;
        RECT -36.900 -77.870 -36.610 -77.820 ;
        RECT -33.570 -77.680 -33.280 -77.630 ;
        RECT -32.210 -77.680 -31.920 -77.620 ;
        RECT -33.570 -77.820 -31.920 -77.680 ;
        RECT -33.570 -77.880 -33.280 -77.820 ;
        RECT -32.210 -77.870 -31.920 -77.820 ;
        RECT -26.790 -77.680 -26.500 -77.620 ;
        RECT -25.400 -77.680 -25.110 -77.620 ;
        RECT -26.790 -77.820 -25.110 -77.680 ;
        RECT -26.790 -77.870 -26.500 -77.820 ;
        RECT -25.400 -77.870 -25.110 -77.820 ;
        RECT -22.070 -77.680 -21.780 -77.630 ;
        RECT -20.710 -77.680 -20.420 -77.620 ;
        RECT -22.070 -77.820 -20.420 -77.680 ;
        RECT -22.070 -77.880 -21.780 -77.820 ;
        RECT -20.710 -77.870 -20.420 -77.820 ;
        RECT -14.970 -77.680 -14.680 -77.620 ;
        RECT -13.580 -77.680 -13.290 -77.620 ;
        RECT -14.970 -77.820 -13.290 -77.680 ;
        RECT -14.970 -77.870 -14.680 -77.820 ;
        RECT -13.580 -77.870 -13.290 -77.820 ;
        RECT -10.250 -77.680 -9.960 -77.630 ;
        RECT -8.890 -77.680 -8.600 -77.620 ;
        RECT -10.250 -77.820 -8.600 -77.680 ;
        RECT -10.250 -77.880 -9.960 -77.820 ;
        RECT -8.890 -77.870 -8.600 -77.820 ;
        RECT -3.160 -77.680 -2.870 -77.620 ;
        RECT -1.770 -77.680 -1.480 -77.620 ;
        RECT -3.160 -77.820 -1.480 -77.680 ;
        RECT -3.160 -77.870 -2.870 -77.820 ;
        RECT -1.770 -77.870 -1.480 -77.820 ;
        RECT 1.560 -77.680 1.850 -77.630 ;
        RECT 2.920 -77.680 3.210 -77.620 ;
        RECT 1.560 -77.820 3.210 -77.680 ;
        RECT 1.560 -77.880 1.850 -77.820 ;
        RECT 2.920 -77.870 3.210 -77.820 ;
        RECT 8.650 -77.680 8.940 -77.620 ;
        RECT 10.040 -77.680 10.330 -77.620 ;
        RECT 8.650 -77.820 10.330 -77.680 ;
        RECT 8.650 -77.870 8.940 -77.820 ;
        RECT 10.040 -77.870 10.330 -77.820 ;
        RECT 13.370 -77.680 13.660 -77.630 ;
        RECT 14.730 -77.680 15.020 -77.620 ;
        RECT 13.370 -77.820 15.020 -77.680 ;
        RECT 13.370 -77.880 13.660 -77.820 ;
        RECT 14.730 -77.870 15.020 -77.820 ;
        RECT 20.470 -77.680 20.760 -77.620 ;
        RECT 21.860 -77.680 22.150 -77.620 ;
        RECT 20.470 -77.820 22.150 -77.680 ;
        RECT 20.470 -77.870 20.760 -77.820 ;
        RECT 21.860 -77.870 22.150 -77.820 ;
        RECT 25.190 -77.680 25.480 -77.630 ;
        RECT 26.550 -77.680 26.840 -77.620 ;
        RECT 25.190 -77.820 26.840 -77.680 ;
        RECT 25.190 -77.880 25.480 -77.820 ;
        RECT 26.550 -77.870 26.840 -77.820 ;
        RECT 32.290 -77.680 32.580 -77.620 ;
        RECT 33.680 -77.680 33.970 -77.620 ;
        RECT 32.290 -77.820 33.970 -77.680 ;
        RECT 32.290 -77.870 32.580 -77.820 ;
        RECT 33.680 -77.870 33.970 -77.820 ;
        RECT 37.010 -77.680 37.300 -77.630 ;
        RECT 38.370 -77.680 38.660 -77.620 ;
        RECT 37.010 -77.820 38.660 -77.680 ;
        RECT 37.010 -77.880 37.300 -77.820 ;
        RECT 38.370 -77.870 38.660 -77.820 ;
        RECT 44.110 -77.680 44.400 -77.620 ;
        RECT 45.500 -77.680 45.790 -77.620 ;
        RECT 44.110 -77.820 45.790 -77.680 ;
        RECT 44.110 -77.870 44.400 -77.820 ;
        RECT 45.500 -77.870 45.790 -77.820 ;
        RECT 48.830 -77.680 49.120 -77.630 ;
        RECT 50.190 -77.680 50.480 -77.620 ;
        RECT 48.830 -77.820 50.480 -77.680 ;
        RECT 48.830 -77.880 49.120 -77.820 ;
        RECT 50.190 -77.870 50.480 -77.820 ;
        RECT 55.930 -77.680 56.220 -77.620 ;
        RECT 57.320 -77.680 57.610 -77.620 ;
        RECT 55.930 -77.820 57.610 -77.680 ;
        RECT 55.930 -77.870 56.220 -77.820 ;
        RECT 57.320 -77.870 57.610 -77.820 ;
        RECT 60.650 -77.680 60.940 -77.630 ;
        RECT 62.010 -77.680 62.300 -77.620 ;
        RECT 60.650 -77.820 62.300 -77.680 ;
        RECT 60.650 -77.880 60.940 -77.820 ;
        RECT 62.010 -77.870 62.300 -77.820 ;
        RECT 67.750 -77.680 68.040 -77.620 ;
        RECT 69.140 -77.680 69.430 -77.620 ;
        RECT 67.750 -77.820 69.430 -77.680 ;
        RECT 67.750 -77.870 68.040 -77.820 ;
        RECT 69.140 -77.870 69.430 -77.820 ;
        RECT 72.470 -77.680 72.760 -77.630 ;
        RECT 73.830 -77.680 74.120 -77.620 ;
        RECT 72.470 -77.820 74.120 -77.680 ;
        RECT 72.470 -77.880 72.760 -77.820 ;
        RECT 73.830 -77.870 74.120 -77.820 ;
        RECT 79.570 -77.680 79.860 -77.620 ;
        RECT 80.960 -77.680 81.250 -77.620 ;
        RECT 79.570 -77.820 81.250 -77.680 ;
        RECT 79.570 -77.870 79.860 -77.820 ;
        RECT 80.960 -77.870 81.250 -77.820 ;
        RECT 84.290 -77.680 84.580 -77.630 ;
        RECT 85.650 -77.680 85.940 -77.620 ;
        RECT 84.290 -77.820 85.940 -77.680 ;
        RECT 84.290 -77.880 84.580 -77.820 ;
        RECT 85.650 -77.870 85.940 -77.820 ;
        RECT 91.410 -77.680 91.700 -77.620 ;
        RECT 92.800 -77.680 93.090 -77.620 ;
        RECT 91.410 -77.820 93.090 -77.680 ;
        RECT 91.410 -77.870 91.700 -77.820 ;
        RECT 92.800 -77.870 93.090 -77.820 ;
        RECT 96.130 -77.680 96.420 -77.630 ;
        RECT 97.490 -77.680 97.780 -77.620 ;
        RECT 96.130 -77.820 97.780 -77.680 ;
        RECT 96.130 -77.880 96.420 -77.820 ;
        RECT 97.490 -77.870 97.780 -77.820 ;
        RECT 103.250 -77.680 103.540 -77.620 ;
        RECT 104.640 -77.680 104.930 -77.620 ;
        RECT 103.250 -77.820 104.930 -77.680 ;
        RECT 103.250 -77.870 103.540 -77.820 ;
        RECT 104.640 -77.870 104.930 -77.820 ;
        RECT 107.970 -77.680 108.260 -77.630 ;
        RECT 109.330 -77.680 109.620 -77.620 ;
        RECT 107.970 -77.820 109.620 -77.680 ;
        RECT 107.970 -77.880 108.260 -77.820 ;
        RECT 109.330 -77.870 109.620 -77.820 ;
        RECT 115.120 -77.680 115.410 -77.620 ;
        RECT 116.510 -77.680 116.800 -77.620 ;
        RECT 115.120 -77.820 116.800 -77.680 ;
        RECT 115.120 -77.870 115.410 -77.820 ;
        RECT 116.510 -77.870 116.800 -77.820 ;
        RECT 119.840 -77.680 120.130 -77.630 ;
        RECT 121.200 -77.680 121.490 -77.620 ;
        RECT 119.840 -77.820 121.490 -77.680 ;
        RECT 119.840 -77.880 120.130 -77.820 ;
        RECT 121.200 -77.870 121.490 -77.820 ;
        RECT 126.990 -77.680 127.280 -77.620 ;
        RECT 128.380 -77.680 128.670 -77.620 ;
        RECT 126.990 -77.820 128.670 -77.680 ;
        RECT 126.990 -77.870 127.280 -77.820 ;
        RECT 128.380 -77.870 128.670 -77.820 ;
        RECT 131.710 -77.680 132.000 -77.630 ;
        RECT 133.070 -77.680 133.360 -77.620 ;
        RECT 131.710 -77.820 133.360 -77.680 ;
        RECT 131.710 -77.880 132.000 -77.820 ;
        RECT 133.070 -77.870 133.360 -77.820 ;
        RECT 136.000 -77.680 136.290 -77.620 ;
        RECT 137.390 -77.680 137.680 -77.620 ;
        RECT 136.000 -77.820 137.680 -77.680 ;
        RECT 136.000 -77.870 136.290 -77.820 ;
        RECT 137.390 -77.870 137.680 -77.820 ;
        RECT 140.720 -77.680 141.010 -77.630 ;
        RECT 142.080 -77.680 142.370 -77.620 ;
        RECT 140.720 -77.820 142.370 -77.680 ;
        RECT 140.720 -77.880 141.010 -77.820 ;
        RECT 142.080 -77.870 142.370 -77.820 ;
        RECT -34.970 -78.420 -34.680 -78.360 ;
        RECT -34.010 -78.420 -33.720 -78.350 ;
        RECT -34.970 -78.560 -33.720 -78.420 ;
        RECT -34.970 -78.610 -34.680 -78.560 ;
        RECT -34.010 -78.600 -33.720 -78.560 ;
        RECT -23.470 -78.420 -23.180 -78.360 ;
        RECT -22.510 -78.420 -22.220 -78.350 ;
        RECT -23.470 -78.560 -22.220 -78.420 ;
        RECT -23.470 -78.610 -23.180 -78.560 ;
        RECT -22.510 -78.600 -22.220 -78.560 ;
        RECT -11.650 -78.420 -11.360 -78.360 ;
        RECT -10.690 -78.420 -10.400 -78.350 ;
        RECT -11.650 -78.560 -10.400 -78.420 ;
        RECT -11.650 -78.610 -11.360 -78.560 ;
        RECT -10.690 -78.600 -10.400 -78.560 ;
        RECT 0.160 -78.420 0.450 -78.360 ;
        RECT 1.120 -78.420 1.410 -78.350 ;
        RECT 0.160 -78.560 1.410 -78.420 ;
        RECT 0.160 -78.610 0.450 -78.560 ;
        RECT 1.120 -78.600 1.410 -78.560 ;
        RECT 11.970 -78.420 12.260 -78.360 ;
        RECT 12.930 -78.420 13.220 -78.350 ;
        RECT 11.970 -78.560 13.220 -78.420 ;
        RECT 11.970 -78.610 12.260 -78.560 ;
        RECT 12.930 -78.600 13.220 -78.560 ;
        RECT 23.790 -78.420 24.080 -78.360 ;
        RECT 24.750 -78.420 25.040 -78.350 ;
        RECT 23.790 -78.560 25.040 -78.420 ;
        RECT 23.790 -78.610 24.080 -78.560 ;
        RECT 24.750 -78.600 25.040 -78.560 ;
        RECT 35.610 -78.420 35.900 -78.360 ;
        RECT 36.570 -78.420 36.860 -78.350 ;
        RECT 35.610 -78.560 36.860 -78.420 ;
        RECT 35.610 -78.610 35.900 -78.560 ;
        RECT 36.570 -78.600 36.860 -78.560 ;
        RECT 47.430 -78.420 47.720 -78.360 ;
        RECT 48.390 -78.420 48.680 -78.350 ;
        RECT 47.430 -78.560 48.680 -78.420 ;
        RECT 47.430 -78.610 47.720 -78.560 ;
        RECT 48.390 -78.600 48.680 -78.560 ;
        RECT 59.250 -78.420 59.540 -78.360 ;
        RECT 60.210 -78.420 60.500 -78.350 ;
        RECT 59.250 -78.560 60.500 -78.420 ;
        RECT 59.250 -78.610 59.540 -78.560 ;
        RECT 60.210 -78.600 60.500 -78.560 ;
        RECT 71.070 -78.420 71.360 -78.360 ;
        RECT 72.030 -78.420 72.320 -78.350 ;
        RECT 71.070 -78.560 72.320 -78.420 ;
        RECT 71.070 -78.610 71.360 -78.560 ;
        RECT 72.030 -78.600 72.320 -78.560 ;
        RECT 82.890 -78.420 83.180 -78.360 ;
        RECT 83.850 -78.420 84.140 -78.350 ;
        RECT 82.890 -78.560 84.140 -78.420 ;
        RECT 82.890 -78.610 83.180 -78.560 ;
        RECT 83.850 -78.600 84.140 -78.560 ;
        RECT 94.730 -78.420 95.020 -78.360 ;
        RECT 95.690 -78.420 95.980 -78.350 ;
        RECT 94.730 -78.560 95.980 -78.420 ;
        RECT 94.730 -78.610 95.020 -78.560 ;
        RECT 95.690 -78.600 95.980 -78.560 ;
        RECT 106.570 -78.420 106.860 -78.360 ;
        RECT 107.530 -78.420 107.820 -78.350 ;
        RECT 106.570 -78.560 107.820 -78.420 ;
        RECT 106.570 -78.610 106.860 -78.560 ;
        RECT 107.530 -78.600 107.820 -78.560 ;
        RECT 118.440 -78.420 118.730 -78.360 ;
        RECT 119.400 -78.420 119.690 -78.350 ;
        RECT 118.440 -78.560 119.690 -78.420 ;
        RECT 118.440 -78.610 118.730 -78.560 ;
        RECT 119.400 -78.600 119.690 -78.560 ;
        RECT 130.310 -78.420 130.600 -78.360 ;
        RECT 131.270 -78.420 131.560 -78.350 ;
        RECT 130.310 -78.560 131.560 -78.420 ;
        RECT 130.310 -78.610 130.600 -78.560 ;
        RECT 131.270 -78.600 131.560 -78.560 ;
        RECT 139.320 -78.420 139.610 -78.360 ;
        RECT 140.280 -78.420 140.570 -78.350 ;
        RECT 139.320 -78.560 140.570 -78.420 ;
        RECT 139.320 -78.610 139.610 -78.560 ;
        RECT 140.280 -78.600 140.570 -78.560 ;
        RECT -36.460 -79.230 -36.170 -79.170 ;
        RECT -35.500 -79.230 -35.210 -79.170 ;
        RECT -36.460 -79.370 -35.210 -79.230 ;
        RECT -36.460 -79.420 -36.170 -79.370 ;
        RECT -35.500 -79.420 -35.210 -79.370 ;
        RECT -24.960 -79.230 -24.670 -79.170 ;
        RECT -24.000 -79.230 -23.710 -79.170 ;
        RECT -24.960 -79.370 -23.710 -79.230 ;
        RECT -24.960 -79.420 -24.670 -79.370 ;
        RECT -24.000 -79.420 -23.710 -79.370 ;
        RECT -13.140 -79.230 -12.850 -79.170 ;
        RECT -12.180 -79.230 -11.890 -79.170 ;
        RECT -13.140 -79.370 -11.890 -79.230 ;
        RECT -13.140 -79.420 -12.850 -79.370 ;
        RECT -12.180 -79.420 -11.890 -79.370 ;
        RECT -1.330 -79.230 -1.040 -79.170 ;
        RECT -0.370 -79.230 -0.080 -79.170 ;
        RECT -1.330 -79.370 -0.080 -79.230 ;
        RECT -1.330 -79.420 -1.040 -79.370 ;
        RECT -0.370 -79.420 -0.080 -79.370 ;
        RECT 10.480 -79.230 10.770 -79.170 ;
        RECT 11.440 -79.230 11.730 -79.170 ;
        RECT 10.480 -79.370 11.730 -79.230 ;
        RECT 10.480 -79.420 10.770 -79.370 ;
        RECT 11.440 -79.420 11.730 -79.370 ;
        RECT 22.300 -79.230 22.590 -79.170 ;
        RECT 23.260 -79.230 23.550 -79.170 ;
        RECT 22.300 -79.370 23.550 -79.230 ;
        RECT 22.300 -79.420 22.590 -79.370 ;
        RECT 23.260 -79.420 23.550 -79.370 ;
        RECT 34.120 -79.230 34.410 -79.170 ;
        RECT 35.080 -79.230 35.370 -79.170 ;
        RECT 34.120 -79.370 35.370 -79.230 ;
        RECT 34.120 -79.420 34.410 -79.370 ;
        RECT 35.080 -79.420 35.370 -79.370 ;
        RECT 45.940 -79.230 46.230 -79.170 ;
        RECT 46.900 -79.230 47.190 -79.170 ;
        RECT 45.940 -79.370 47.190 -79.230 ;
        RECT 45.940 -79.420 46.230 -79.370 ;
        RECT 46.900 -79.420 47.190 -79.370 ;
        RECT 57.760 -79.230 58.050 -79.170 ;
        RECT 58.720 -79.230 59.010 -79.170 ;
        RECT 57.760 -79.370 59.010 -79.230 ;
        RECT 57.760 -79.420 58.050 -79.370 ;
        RECT 58.720 -79.420 59.010 -79.370 ;
        RECT 69.580 -79.230 69.870 -79.170 ;
        RECT 70.540 -79.230 70.830 -79.170 ;
        RECT 69.580 -79.370 70.830 -79.230 ;
        RECT 69.580 -79.420 69.870 -79.370 ;
        RECT 70.540 -79.420 70.830 -79.370 ;
        RECT 81.400 -79.230 81.690 -79.170 ;
        RECT 82.360 -79.230 82.650 -79.170 ;
        RECT 81.400 -79.370 82.650 -79.230 ;
        RECT 81.400 -79.420 81.690 -79.370 ;
        RECT 82.360 -79.420 82.650 -79.370 ;
        RECT 93.240 -79.230 93.530 -79.170 ;
        RECT 94.200 -79.230 94.490 -79.170 ;
        RECT 93.240 -79.370 94.490 -79.230 ;
        RECT 93.240 -79.420 93.530 -79.370 ;
        RECT 94.200 -79.420 94.490 -79.370 ;
        RECT 105.080 -79.230 105.370 -79.170 ;
        RECT 106.040 -79.230 106.330 -79.170 ;
        RECT 105.080 -79.370 106.330 -79.230 ;
        RECT 105.080 -79.420 105.370 -79.370 ;
        RECT 106.040 -79.420 106.330 -79.370 ;
        RECT 116.950 -79.230 117.240 -79.170 ;
        RECT 117.910 -79.230 118.200 -79.170 ;
        RECT 116.950 -79.370 118.200 -79.230 ;
        RECT 116.950 -79.420 117.240 -79.370 ;
        RECT 117.910 -79.420 118.200 -79.370 ;
        RECT 128.820 -79.230 129.110 -79.170 ;
        RECT 129.780 -79.230 130.070 -79.170 ;
        RECT 128.820 -79.370 130.070 -79.230 ;
        RECT 128.820 -79.420 129.110 -79.370 ;
        RECT 129.780 -79.420 130.070 -79.370 ;
        RECT 137.830 -79.230 138.120 -79.170 ;
        RECT 138.790 -79.230 139.080 -79.170 ;
        RECT 137.830 -79.370 139.080 -79.230 ;
        RECT 137.830 -79.420 138.120 -79.370 ;
        RECT 138.790 -79.420 139.080 -79.370 ;
        RECT -37.940 -79.900 -37.650 -79.850 ;
        RECT -36.460 -79.900 -36.170 -79.880 ;
        RECT -37.940 -80.040 -36.170 -79.900 ;
        RECT -37.940 -80.100 -37.650 -80.040 ;
        RECT -36.460 -80.130 -36.170 -80.040 ;
        RECT -34.010 -79.930 -33.720 -79.890 ;
        RECT -32.560 -79.930 -32.270 -79.860 ;
        RECT -34.010 -80.070 -32.270 -79.930 ;
        RECT -34.010 -80.140 -33.720 -80.070 ;
        RECT -32.560 -80.110 -32.270 -80.070 ;
        RECT -26.440 -79.900 -26.150 -79.850 ;
        RECT -24.960 -79.900 -24.670 -79.880 ;
        RECT -26.440 -80.040 -24.670 -79.900 ;
        RECT -26.440 -80.100 -26.150 -80.040 ;
        RECT -24.960 -80.130 -24.670 -80.040 ;
        RECT -22.510 -79.930 -22.220 -79.890 ;
        RECT -21.060 -79.930 -20.770 -79.860 ;
        RECT -22.510 -80.070 -20.770 -79.930 ;
        RECT -22.510 -80.140 -22.220 -80.070 ;
        RECT -21.060 -80.110 -20.770 -80.070 ;
        RECT -14.620 -79.900 -14.330 -79.850 ;
        RECT -13.140 -79.900 -12.850 -79.880 ;
        RECT -14.620 -80.040 -12.850 -79.900 ;
        RECT -14.620 -80.100 -14.330 -80.040 ;
        RECT -13.140 -80.130 -12.850 -80.040 ;
        RECT -10.690 -79.930 -10.400 -79.890 ;
        RECT -9.240 -79.930 -8.950 -79.860 ;
        RECT -10.690 -80.070 -8.950 -79.930 ;
        RECT -10.690 -80.140 -10.400 -80.070 ;
        RECT -9.240 -80.110 -8.950 -80.070 ;
        RECT -2.810 -79.900 -2.520 -79.850 ;
        RECT -1.330 -79.900 -1.040 -79.880 ;
        RECT -2.810 -80.040 -1.040 -79.900 ;
        RECT -2.810 -80.100 -2.520 -80.040 ;
        RECT -1.330 -80.130 -1.040 -80.040 ;
        RECT 1.120 -79.930 1.410 -79.890 ;
        RECT 2.570 -79.930 2.860 -79.860 ;
        RECT 1.120 -80.070 2.860 -79.930 ;
        RECT 1.120 -80.140 1.410 -80.070 ;
        RECT 2.570 -80.110 2.860 -80.070 ;
        RECT 9.000 -79.900 9.290 -79.850 ;
        RECT 10.480 -79.900 10.770 -79.880 ;
        RECT 9.000 -80.040 10.770 -79.900 ;
        RECT 9.000 -80.100 9.290 -80.040 ;
        RECT 10.480 -80.130 10.770 -80.040 ;
        RECT 12.930 -79.930 13.220 -79.890 ;
        RECT 14.380 -79.930 14.670 -79.860 ;
        RECT 12.930 -80.070 14.670 -79.930 ;
        RECT 12.930 -80.140 13.220 -80.070 ;
        RECT 14.380 -80.110 14.670 -80.070 ;
        RECT 20.820 -79.900 21.110 -79.850 ;
        RECT 22.300 -79.900 22.590 -79.880 ;
        RECT 20.820 -80.040 22.590 -79.900 ;
        RECT 20.820 -80.100 21.110 -80.040 ;
        RECT 22.300 -80.130 22.590 -80.040 ;
        RECT 24.750 -79.930 25.040 -79.890 ;
        RECT 26.200 -79.930 26.490 -79.860 ;
        RECT 24.750 -80.070 26.490 -79.930 ;
        RECT 24.750 -80.140 25.040 -80.070 ;
        RECT 26.200 -80.110 26.490 -80.070 ;
        RECT 32.640 -79.900 32.930 -79.850 ;
        RECT 34.120 -79.900 34.410 -79.880 ;
        RECT 32.640 -80.040 34.410 -79.900 ;
        RECT 32.640 -80.100 32.930 -80.040 ;
        RECT 34.120 -80.130 34.410 -80.040 ;
        RECT 36.570 -79.930 36.860 -79.890 ;
        RECT 38.020 -79.930 38.310 -79.860 ;
        RECT 36.570 -80.070 38.310 -79.930 ;
        RECT 36.570 -80.140 36.860 -80.070 ;
        RECT 38.020 -80.110 38.310 -80.070 ;
        RECT 44.460 -79.900 44.750 -79.850 ;
        RECT 45.940 -79.900 46.230 -79.880 ;
        RECT 44.460 -80.040 46.230 -79.900 ;
        RECT 44.460 -80.100 44.750 -80.040 ;
        RECT 45.940 -80.130 46.230 -80.040 ;
        RECT 48.390 -79.930 48.680 -79.890 ;
        RECT 49.840 -79.930 50.130 -79.860 ;
        RECT 48.390 -80.070 50.130 -79.930 ;
        RECT 48.390 -80.140 48.680 -80.070 ;
        RECT 49.840 -80.110 50.130 -80.070 ;
        RECT 56.280 -79.900 56.570 -79.850 ;
        RECT 57.760 -79.900 58.050 -79.880 ;
        RECT 56.280 -80.040 58.050 -79.900 ;
        RECT 56.280 -80.100 56.570 -80.040 ;
        RECT 57.760 -80.130 58.050 -80.040 ;
        RECT 60.210 -79.930 60.500 -79.890 ;
        RECT 61.660 -79.930 61.950 -79.860 ;
        RECT 60.210 -80.070 61.950 -79.930 ;
        RECT 60.210 -80.140 60.500 -80.070 ;
        RECT 61.660 -80.110 61.950 -80.070 ;
        RECT 68.100 -79.900 68.390 -79.850 ;
        RECT 69.580 -79.900 69.870 -79.880 ;
        RECT 68.100 -80.040 69.870 -79.900 ;
        RECT 68.100 -80.100 68.390 -80.040 ;
        RECT 69.580 -80.130 69.870 -80.040 ;
        RECT 72.030 -79.930 72.320 -79.890 ;
        RECT 73.480 -79.930 73.770 -79.860 ;
        RECT 72.030 -80.070 73.770 -79.930 ;
        RECT 72.030 -80.140 72.320 -80.070 ;
        RECT 73.480 -80.110 73.770 -80.070 ;
        RECT 79.920 -79.900 80.210 -79.850 ;
        RECT 81.400 -79.900 81.690 -79.880 ;
        RECT 79.920 -80.040 81.690 -79.900 ;
        RECT 79.920 -80.100 80.210 -80.040 ;
        RECT 81.400 -80.130 81.690 -80.040 ;
        RECT 83.850 -79.930 84.140 -79.890 ;
        RECT 85.300 -79.930 85.590 -79.860 ;
        RECT 83.850 -80.070 85.590 -79.930 ;
        RECT 83.850 -80.140 84.140 -80.070 ;
        RECT 85.300 -80.110 85.590 -80.070 ;
        RECT 91.760 -79.900 92.050 -79.850 ;
        RECT 93.240 -79.900 93.530 -79.880 ;
        RECT 91.760 -80.040 93.530 -79.900 ;
        RECT 91.760 -80.100 92.050 -80.040 ;
        RECT 93.240 -80.130 93.530 -80.040 ;
        RECT 95.690 -79.930 95.980 -79.890 ;
        RECT 97.140 -79.930 97.430 -79.860 ;
        RECT 95.690 -80.070 97.430 -79.930 ;
        RECT 95.690 -80.140 95.980 -80.070 ;
        RECT 97.140 -80.110 97.430 -80.070 ;
        RECT 103.600 -79.900 103.890 -79.850 ;
        RECT 105.080 -79.900 105.370 -79.880 ;
        RECT 103.600 -80.040 105.370 -79.900 ;
        RECT 103.600 -80.100 103.890 -80.040 ;
        RECT 105.080 -80.130 105.370 -80.040 ;
        RECT 107.530 -79.930 107.820 -79.890 ;
        RECT 108.980 -79.930 109.270 -79.860 ;
        RECT 107.530 -80.070 109.270 -79.930 ;
        RECT 107.530 -80.140 107.820 -80.070 ;
        RECT 108.980 -80.110 109.270 -80.070 ;
        RECT 115.470 -79.900 115.760 -79.850 ;
        RECT 116.950 -79.900 117.240 -79.880 ;
        RECT 115.470 -80.040 117.240 -79.900 ;
        RECT 115.470 -80.100 115.760 -80.040 ;
        RECT 116.950 -80.130 117.240 -80.040 ;
        RECT 119.400 -79.930 119.690 -79.890 ;
        RECT 120.850 -79.930 121.140 -79.860 ;
        RECT 119.400 -80.070 121.140 -79.930 ;
        RECT 119.400 -80.140 119.690 -80.070 ;
        RECT 120.850 -80.110 121.140 -80.070 ;
        RECT 127.340 -79.900 127.630 -79.850 ;
        RECT 128.820 -79.900 129.110 -79.880 ;
        RECT 127.340 -80.040 129.110 -79.900 ;
        RECT 127.340 -80.100 127.630 -80.040 ;
        RECT 128.820 -80.130 129.110 -80.040 ;
        RECT 131.270 -79.930 131.560 -79.890 ;
        RECT 132.720 -79.930 133.010 -79.860 ;
        RECT 131.270 -80.070 133.010 -79.930 ;
        RECT 131.270 -80.140 131.560 -80.070 ;
        RECT 132.720 -80.110 133.010 -80.070 ;
        RECT 136.350 -79.900 136.640 -79.850 ;
        RECT 137.830 -79.900 138.120 -79.880 ;
        RECT 136.350 -80.040 138.120 -79.900 ;
        RECT 136.350 -80.100 136.640 -80.040 ;
        RECT 137.830 -80.130 138.120 -80.040 ;
        RECT 140.280 -79.930 140.570 -79.890 ;
        RECT 141.730 -79.930 142.020 -79.860 ;
        RECT 140.280 -80.070 142.020 -79.930 ;
        RECT 140.280 -80.140 140.570 -80.070 ;
        RECT 141.730 -80.110 142.020 -80.070 ;
        RECT -41.230 -80.530 -40.910 -80.470 ;
        RECT -37.860 -80.520 -37.570 -80.490 ;
        RECT -37.900 -80.530 -37.570 -80.520 ;
        RECT -32.640 -80.500 -32.350 -80.470 ;
        RECT -32.640 -80.530 -32.310 -80.500 ;
        RECT -26.360 -80.520 -26.070 -80.490 ;
        RECT -26.400 -80.530 -26.070 -80.520 ;
        RECT -21.140 -80.500 -20.850 -80.470 ;
        RECT -21.140 -80.530 -20.810 -80.500 ;
        RECT -14.540 -80.520 -14.250 -80.490 ;
        RECT -14.580 -80.530 -14.250 -80.520 ;
        RECT -9.320 -80.500 -9.030 -80.470 ;
        RECT -9.320 -80.530 -8.990 -80.500 ;
        RECT -2.730 -80.520 -2.440 -80.490 ;
        RECT -2.770 -80.530 -2.440 -80.520 ;
        RECT 2.490 -80.500 2.780 -80.470 ;
        RECT 2.490 -80.530 2.820 -80.500 ;
        RECT 9.080 -80.520 9.370 -80.490 ;
        RECT 9.040 -80.530 9.370 -80.520 ;
        RECT 14.300 -80.500 14.590 -80.470 ;
        RECT 14.300 -80.530 14.630 -80.500 ;
        RECT 20.900 -80.520 21.190 -80.490 ;
        RECT 20.860 -80.530 21.190 -80.520 ;
        RECT 26.120 -80.500 26.410 -80.470 ;
        RECT 26.120 -80.530 26.450 -80.500 ;
        RECT 32.720 -80.520 33.010 -80.490 ;
        RECT 32.680 -80.530 33.010 -80.520 ;
        RECT 37.940 -80.500 38.230 -80.470 ;
        RECT 37.940 -80.530 38.270 -80.500 ;
        RECT 44.540 -80.520 44.830 -80.490 ;
        RECT 44.500 -80.530 44.830 -80.520 ;
        RECT 49.760 -80.500 50.050 -80.470 ;
        RECT 49.760 -80.530 50.090 -80.500 ;
        RECT 56.360 -80.520 56.650 -80.490 ;
        RECT 56.320 -80.530 56.650 -80.520 ;
        RECT 61.580 -80.500 61.870 -80.470 ;
        RECT 61.580 -80.530 61.910 -80.500 ;
        RECT 68.180 -80.520 68.470 -80.490 ;
        RECT 68.140 -80.530 68.470 -80.520 ;
        RECT 73.400 -80.500 73.690 -80.470 ;
        RECT 73.400 -80.530 73.730 -80.500 ;
        RECT 80.000 -80.520 80.290 -80.490 ;
        RECT 79.960 -80.530 80.290 -80.520 ;
        RECT 85.220 -80.500 85.510 -80.470 ;
        RECT 85.220 -80.530 85.550 -80.500 ;
        RECT 91.840 -80.520 92.130 -80.490 ;
        RECT 91.800 -80.530 92.130 -80.520 ;
        RECT 97.060 -80.500 97.350 -80.470 ;
        RECT 97.060 -80.530 97.390 -80.500 ;
        RECT 103.680 -80.520 103.970 -80.490 ;
        RECT 103.640 -80.530 103.970 -80.520 ;
        RECT 108.900 -80.500 109.190 -80.470 ;
        RECT 108.900 -80.530 109.230 -80.500 ;
        RECT 115.550 -80.520 115.840 -80.490 ;
        RECT 115.510 -80.530 115.840 -80.520 ;
        RECT 120.770 -80.500 121.060 -80.470 ;
        RECT 120.770 -80.530 121.100 -80.500 ;
        RECT 127.420 -80.520 127.710 -80.490 ;
        RECT 127.380 -80.530 127.710 -80.520 ;
        RECT 132.640 -80.500 132.930 -80.470 ;
        RECT 132.640 -80.530 132.970 -80.500 ;
        RECT 136.430 -80.520 136.720 -80.490 ;
        RECT 136.390 -80.530 136.720 -80.520 ;
        RECT 141.650 -80.500 141.940 -80.470 ;
        RECT 141.650 -80.530 141.980 -80.500 ;
        RECT -41.230 -80.670 142.470 -80.530 ;
        RECT -41.230 -80.730 -40.910 -80.670 ;
        RECT -37.900 -80.700 -37.570 -80.670 ;
        RECT -37.860 -80.730 -37.570 -80.700 ;
        RECT -32.640 -80.680 -32.310 -80.670 ;
        RECT -32.640 -80.710 -32.350 -80.680 ;
        RECT -26.400 -80.700 -26.070 -80.670 ;
        RECT -26.360 -80.730 -26.070 -80.700 ;
        RECT -21.140 -80.680 -20.810 -80.670 ;
        RECT -21.140 -80.710 -20.850 -80.680 ;
        RECT -14.580 -80.700 -14.250 -80.670 ;
        RECT -14.540 -80.730 -14.250 -80.700 ;
        RECT -9.320 -80.680 -8.990 -80.670 ;
        RECT -9.320 -80.710 -9.030 -80.680 ;
        RECT -2.770 -80.700 -2.440 -80.670 ;
        RECT -2.730 -80.730 -2.440 -80.700 ;
        RECT 2.490 -80.680 2.820 -80.670 ;
        RECT 2.490 -80.710 2.780 -80.680 ;
        RECT 9.040 -80.700 9.370 -80.670 ;
        RECT 9.080 -80.730 9.370 -80.700 ;
        RECT 14.300 -80.680 14.630 -80.670 ;
        RECT 14.300 -80.710 14.590 -80.680 ;
        RECT 20.860 -80.700 21.190 -80.670 ;
        RECT 20.900 -80.730 21.190 -80.700 ;
        RECT 26.120 -80.680 26.450 -80.670 ;
        RECT 26.120 -80.710 26.410 -80.680 ;
        RECT 32.680 -80.700 33.010 -80.670 ;
        RECT 32.720 -80.730 33.010 -80.700 ;
        RECT 37.940 -80.680 38.270 -80.670 ;
        RECT 37.940 -80.710 38.230 -80.680 ;
        RECT 44.500 -80.700 44.830 -80.670 ;
        RECT 44.540 -80.730 44.830 -80.700 ;
        RECT 49.760 -80.680 50.090 -80.670 ;
        RECT 49.760 -80.710 50.050 -80.680 ;
        RECT 56.320 -80.700 56.650 -80.670 ;
        RECT 56.360 -80.730 56.650 -80.700 ;
        RECT 61.580 -80.680 61.910 -80.670 ;
        RECT 61.580 -80.710 61.870 -80.680 ;
        RECT 68.140 -80.700 68.470 -80.670 ;
        RECT 68.180 -80.730 68.470 -80.700 ;
        RECT 73.400 -80.680 73.730 -80.670 ;
        RECT 73.400 -80.710 73.690 -80.680 ;
        RECT 79.960 -80.700 80.290 -80.670 ;
        RECT 80.000 -80.730 80.290 -80.700 ;
        RECT 85.220 -80.680 85.550 -80.670 ;
        RECT 85.220 -80.710 85.510 -80.680 ;
        RECT 91.800 -80.700 92.130 -80.670 ;
        RECT 91.840 -80.730 92.130 -80.700 ;
        RECT 97.060 -80.680 97.390 -80.670 ;
        RECT 97.060 -80.710 97.350 -80.680 ;
        RECT 103.640 -80.700 103.970 -80.670 ;
        RECT 103.680 -80.730 103.970 -80.700 ;
        RECT 108.900 -80.680 109.230 -80.670 ;
        RECT 108.900 -80.710 109.190 -80.680 ;
        RECT 115.510 -80.700 115.840 -80.670 ;
        RECT 115.550 -80.730 115.840 -80.700 ;
        RECT 120.770 -80.680 121.100 -80.670 ;
        RECT 120.770 -80.710 121.060 -80.680 ;
        RECT 127.380 -80.700 127.710 -80.670 ;
        RECT 127.420 -80.730 127.710 -80.700 ;
        RECT 132.640 -80.680 132.970 -80.670 ;
        RECT 132.640 -80.710 132.930 -80.680 ;
        RECT 136.390 -80.700 136.720 -80.670 ;
        RECT 136.430 -80.730 136.720 -80.700 ;
        RECT 141.650 -80.680 141.980 -80.670 ;
        RECT 141.650 -80.710 141.940 -80.680 ;
        RECT -40.570 -80.930 -40.250 -80.870 ;
        RECT -36.790 -80.930 -36.460 -80.880 ;
        RECT -33.720 -80.930 -33.390 -80.890 ;
        RECT -25.290 -80.930 -24.960 -80.880 ;
        RECT -22.220 -80.930 -21.890 -80.890 ;
        RECT -13.470 -80.930 -13.140 -80.880 ;
        RECT -10.400 -80.930 -10.070 -80.890 ;
        RECT -1.660 -80.930 -1.330 -80.880 ;
        RECT 1.410 -80.930 1.740 -80.890 ;
        RECT 10.150 -80.930 10.480 -80.880 ;
        RECT 13.220 -80.930 13.550 -80.890 ;
        RECT 21.970 -80.930 22.300 -80.880 ;
        RECT 25.040 -80.930 25.370 -80.890 ;
        RECT 33.790 -80.930 34.120 -80.880 ;
        RECT 36.860 -80.930 37.190 -80.890 ;
        RECT 45.610 -80.930 45.940 -80.880 ;
        RECT 48.680 -80.930 49.010 -80.890 ;
        RECT 57.430 -80.930 57.760 -80.880 ;
        RECT 60.500 -80.930 60.830 -80.890 ;
        RECT 69.250 -80.930 69.580 -80.880 ;
        RECT 72.320 -80.930 72.650 -80.890 ;
        RECT 81.070 -80.930 81.400 -80.880 ;
        RECT 84.140 -80.930 84.470 -80.890 ;
        RECT 92.910 -80.930 93.240 -80.880 ;
        RECT 95.980 -80.930 96.310 -80.890 ;
        RECT 104.750 -80.930 105.080 -80.880 ;
        RECT 107.820 -80.930 108.150 -80.890 ;
        RECT 116.620 -80.930 116.950 -80.880 ;
        RECT 119.690 -80.930 120.020 -80.890 ;
        RECT 128.490 -80.930 128.820 -80.880 ;
        RECT 131.560 -80.930 131.890 -80.890 ;
        RECT 137.500 -80.930 137.830 -80.880 ;
        RECT 140.570 -80.930 140.900 -80.890 ;
        RECT -40.570 -81.070 142.470 -80.930 ;
        RECT -40.570 -81.130 -40.250 -81.070 ;
        RECT -36.790 -81.120 -36.460 -81.070 ;
        RECT -33.720 -81.130 -33.390 -81.070 ;
        RECT -25.290 -81.120 -24.960 -81.070 ;
        RECT -22.220 -81.130 -21.890 -81.070 ;
        RECT -13.470 -81.120 -13.140 -81.070 ;
        RECT -10.400 -81.130 -10.070 -81.070 ;
        RECT -1.660 -81.120 -1.330 -81.070 ;
        RECT 1.410 -81.130 1.740 -81.070 ;
        RECT 10.150 -81.120 10.480 -81.070 ;
        RECT 13.220 -81.130 13.550 -81.070 ;
        RECT 21.970 -81.120 22.300 -81.070 ;
        RECT 25.040 -81.130 25.370 -81.070 ;
        RECT 33.790 -81.120 34.120 -81.070 ;
        RECT 36.860 -81.130 37.190 -81.070 ;
        RECT 45.610 -81.120 45.940 -81.070 ;
        RECT 48.680 -81.130 49.010 -81.070 ;
        RECT 57.430 -81.120 57.760 -81.070 ;
        RECT 60.500 -81.130 60.830 -81.070 ;
        RECT 69.250 -81.120 69.580 -81.070 ;
        RECT 72.320 -81.130 72.650 -81.070 ;
        RECT 81.070 -81.120 81.400 -81.070 ;
        RECT 84.140 -81.130 84.470 -81.070 ;
        RECT 92.910 -81.120 93.240 -81.070 ;
        RECT 95.980 -81.130 96.310 -81.070 ;
        RECT 104.750 -81.120 105.080 -81.070 ;
        RECT 107.820 -81.130 108.150 -81.070 ;
        RECT 116.620 -81.120 116.950 -81.070 ;
        RECT 119.690 -81.130 120.020 -81.070 ;
        RECT 128.490 -81.120 128.820 -81.070 ;
        RECT 131.560 -81.130 131.890 -81.070 ;
        RECT 137.500 -81.120 137.830 -81.070 ;
        RECT 140.570 -81.130 140.900 -81.070 ;
        RECT -36.460 -81.360 -36.230 -81.290 ;
        RECT -30.290 -81.360 -29.970 -81.300 ;
        RECT -36.460 -81.500 -29.970 -81.360 ;
        RECT -36.460 -81.580 -36.230 -81.500 ;
        RECT -30.290 -81.560 -29.970 -81.500 ;
        RECT -25.140 -81.360 -24.850 -81.290 ;
        RECT -18.730 -81.360 -18.410 -81.300 ;
        RECT -25.140 -81.500 -18.410 -81.360 ;
        RECT -25.140 -81.580 -24.850 -81.500 ;
        RECT -18.730 -81.560 -18.410 -81.500 ;
        RECT -13.390 -81.360 -13.100 -81.290 ;
        RECT -7.040 -81.360 -6.720 -81.300 ;
        RECT -13.390 -81.500 -6.720 -81.360 ;
        RECT -13.390 -81.580 -13.100 -81.500 ;
        RECT -7.040 -81.560 -6.720 -81.500 ;
        RECT -1.570 -81.360 -1.280 -81.290 ;
        RECT 4.870 -81.360 5.190 -81.300 ;
        RECT -1.570 -81.500 5.190 -81.360 ;
        RECT -1.570 -81.580 -1.280 -81.500 ;
        RECT 4.870 -81.560 5.190 -81.500 ;
        RECT 10.250 -81.360 10.540 -81.290 ;
        RECT 16.640 -81.360 16.960 -81.300 ;
        RECT 10.250 -81.500 16.960 -81.360 ;
        RECT 10.250 -81.580 10.540 -81.500 ;
        RECT 16.640 -81.560 16.960 -81.500 ;
        RECT 22.070 -81.360 22.360 -81.290 ;
        RECT 28.410 -81.360 28.730 -81.300 ;
        RECT 22.070 -81.500 28.730 -81.360 ;
        RECT 22.070 -81.580 22.360 -81.500 ;
        RECT 28.410 -81.560 28.730 -81.500 ;
        RECT 34.010 -81.360 34.300 -81.290 ;
        RECT 40.230 -81.360 40.550 -81.300 ;
        RECT 34.010 -81.500 40.550 -81.360 ;
        RECT 34.010 -81.580 34.300 -81.500 ;
        RECT 40.230 -81.560 40.550 -81.500 ;
        RECT 45.780 -81.360 46.070 -81.290 ;
        RECT 52.090 -81.360 52.410 -81.300 ;
        RECT 45.780 -81.500 52.410 -81.360 ;
        RECT 45.780 -81.580 46.070 -81.500 ;
        RECT 52.090 -81.560 52.410 -81.500 ;
        RECT 57.610 -81.360 57.900 -81.290 ;
        RECT 63.880 -81.360 64.200 -81.300 ;
        RECT 57.610 -81.500 64.200 -81.360 ;
        RECT 57.610 -81.580 57.900 -81.500 ;
        RECT 63.880 -81.560 64.200 -81.500 ;
        RECT 69.340 -81.360 69.630 -81.290 ;
        RECT 75.760 -81.360 76.080 -81.300 ;
        RECT 69.340 -81.500 76.080 -81.360 ;
        RECT 69.340 -81.580 69.630 -81.500 ;
        RECT 75.760 -81.560 76.080 -81.500 ;
        RECT 81.170 -81.360 81.460 -81.290 ;
        RECT 87.490 -81.360 87.810 -81.300 ;
        RECT 81.170 -81.500 87.810 -81.360 ;
        RECT 81.170 -81.580 81.460 -81.500 ;
        RECT 87.490 -81.560 87.810 -81.500 ;
        RECT 93.000 -81.360 93.290 -81.290 ;
        RECT 99.310 -81.360 99.630 -81.300 ;
        RECT 93.000 -81.500 99.630 -81.360 ;
        RECT 93.000 -81.580 93.290 -81.500 ;
        RECT 99.310 -81.560 99.630 -81.500 ;
        RECT 104.780 -81.360 105.070 -81.290 ;
        RECT 111.200 -81.360 111.520 -81.300 ;
        RECT 104.780 -81.500 111.520 -81.360 ;
        RECT 104.780 -81.580 105.070 -81.500 ;
        RECT 111.200 -81.560 111.520 -81.500 ;
        RECT 116.720 -81.360 117.010 -81.290 ;
        RECT 123.150 -81.360 123.470 -81.300 ;
        RECT 116.720 -81.500 123.470 -81.360 ;
        RECT 116.720 -81.580 117.010 -81.500 ;
        RECT 123.150 -81.560 123.470 -81.500 ;
        RECT 128.670 -81.360 128.960 -81.290 ;
        RECT 134.910 -81.360 135.230 -81.300 ;
        RECT 128.670 -81.500 135.230 -81.360 ;
        RECT 128.670 -81.580 128.960 -81.500 ;
        RECT 134.910 -81.560 135.230 -81.500 ;
        RECT 137.720 -81.360 138.010 -81.290 ;
        RECT 143.950 -81.360 144.270 -81.300 ;
        RECT 137.720 -81.500 144.270 -81.360 ;
        RECT 137.720 -81.580 138.010 -81.500 ;
        RECT 143.950 -81.560 144.270 -81.500 ;
        RECT -37.000 -83.600 -36.750 -83.490 ;
        RECT -35.250 -83.600 -34.930 -83.510 ;
        RECT -37.000 -83.610 -34.930 -83.600 ;
        RECT -33.460 -83.610 -33.210 -83.520 ;
        RECT -32.400 -83.610 -32.110 -83.560 ;
        RECT -37.000 -83.740 -32.110 -83.610 ;
        RECT -37.000 -83.850 -36.750 -83.740 ;
        RECT -35.250 -83.750 -32.110 -83.740 ;
        RECT -35.250 -83.830 -34.930 -83.750 ;
        RECT -33.460 -83.840 -33.210 -83.750 ;
        RECT -32.400 -83.790 -32.110 -83.750 ;
        RECT -25.500 -83.600 -25.250 -83.490 ;
        RECT -23.750 -83.600 -23.430 -83.510 ;
        RECT -25.500 -83.610 -23.430 -83.600 ;
        RECT -21.960 -83.610 -21.710 -83.520 ;
        RECT -20.900 -83.610 -20.610 -83.560 ;
        RECT -25.500 -83.740 -20.610 -83.610 ;
        RECT -25.500 -83.850 -25.250 -83.740 ;
        RECT -23.750 -83.750 -20.610 -83.740 ;
        RECT -23.750 -83.830 -23.430 -83.750 ;
        RECT -21.960 -83.840 -21.710 -83.750 ;
        RECT -20.900 -83.790 -20.610 -83.750 ;
        RECT -13.680 -83.600 -13.430 -83.490 ;
        RECT -11.930 -83.600 -11.610 -83.510 ;
        RECT -13.680 -83.610 -11.610 -83.600 ;
        RECT -10.140 -83.610 -9.890 -83.520 ;
        RECT -9.080 -83.610 -8.790 -83.560 ;
        RECT -13.680 -83.740 -8.790 -83.610 ;
        RECT -13.680 -83.850 -13.430 -83.740 ;
        RECT -11.930 -83.750 -8.790 -83.740 ;
        RECT -11.930 -83.830 -11.610 -83.750 ;
        RECT -10.140 -83.840 -9.890 -83.750 ;
        RECT -9.080 -83.790 -8.790 -83.750 ;
        RECT -1.870 -83.600 -1.620 -83.490 ;
        RECT -0.120 -83.600 0.200 -83.510 ;
        RECT -1.870 -83.610 0.200 -83.600 ;
        RECT 1.670 -83.610 1.920 -83.520 ;
        RECT 2.730 -83.610 3.020 -83.560 ;
        RECT -1.870 -83.740 3.020 -83.610 ;
        RECT -1.870 -83.850 -1.620 -83.740 ;
        RECT -0.120 -83.750 3.020 -83.740 ;
        RECT -0.120 -83.830 0.200 -83.750 ;
        RECT 1.670 -83.840 1.920 -83.750 ;
        RECT 2.730 -83.790 3.020 -83.750 ;
        RECT 9.940 -83.600 10.190 -83.490 ;
        RECT 11.690 -83.600 12.010 -83.510 ;
        RECT 9.940 -83.610 12.010 -83.600 ;
        RECT 13.480 -83.610 13.730 -83.520 ;
        RECT 14.540 -83.610 14.830 -83.560 ;
        RECT 9.940 -83.740 14.830 -83.610 ;
        RECT 9.940 -83.850 10.190 -83.740 ;
        RECT 11.690 -83.750 14.830 -83.740 ;
        RECT 11.690 -83.830 12.010 -83.750 ;
        RECT 13.480 -83.840 13.730 -83.750 ;
        RECT 14.540 -83.790 14.830 -83.750 ;
        RECT 21.760 -83.600 22.010 -83.490 ;
        RECT 23.510 -83.600 23.830 -83.510 ;
        RECT 21.760 -83.610 23.830 -83.600 ;
        RECT 25.300 -83.610 25.550 -83.520 ;
        RECT 26.360 -83.610 26.650 -83.560 ;
        RECT 21.760 -83.740 26.650 -83.610 ;
        RECT 21.760 -83.850 22.010 -83.740 ;
        RECT 23.510 -83.750 26.650 -83.740 ;
        RECT 23.510 -83.830 23.830 -83.750 ;
        RECT 25.300 -83.840 25.550 -83.750 ;
        RECT 26.360 -83.790 26.650 -83.750 ;
        RECT 33.580 -83.600 33.830 -83.490 ;
        RECT 35.330 -83.600 35.650 -83.510 ;
        RECT 33.580 -83.610 35.650 -83.600 ;
        RECT 37.120 -83.610 37.370 -83.520 ;
        RECT 38.180 -83.610 38.470 -83.560 ;
        RECT 33.580 -83.740 38.470 -83.610 ;
        RECT 33.580 -83.850 33.830 -83.740 ;
        RECT 35.330 -83.750 38.470 -83.740 ;
        RECT 35.330 -83.830 35.650 -83.750 ;
        RECT 37.120 -83.840 37.370 -83.750 ;
        RECT 38.180 -83.790 38.470 -83.750 ;
        RECT 45.400 -83.600 45.650 -83.490 ;
        RECT 47.150 -83.600 47.470 -83.510 ;
        RECT 45.400 -83.610 47.470 -83.600 ;
        RECT 48.940 -83.610 49.190 -83.520 ;
        RECT 50.000 -83.610 50.290 -83.560 ;
        RECT 45.400 -83.740 50.290 -83.610 ;
        RECT 45.400 -83.850 45.650 -83.740 ;
        RECT 47.150 -83.750 50.290 -83.740 ;
        RECT 47.150 -83.830 47.470 -83.750 ;
        RECT 48.940 -83.840 49.190 -83.750 ;
        RECT 50.000 -83.790 50.290 -83.750 ;
        RECT 57.220 -83.600 57.470 -83.490 ;
        RECT 58.970 -83.600 59.290 -83.510 ;
        RECT 57.220 -83.610 59.290 -83.600 ;
        RECT 60.760 -83.610 61.010 -83.520 ;
        RECT 61.820 -83.610 62.110 -83.560 ;
        RECT 57.220 -83.740 62.110 -83.610 ;
        RECT 57.220 -83.850 57.470 -83.740 ;
        RECT 58.970 -83.750 62.110 -83.740 ;
        RECT 58.970 -83.830 59.290 -83.750 ;
        RECT 60.760 -83.840 61.010 -83.750 ;
        RECT 61.820 -83.790 62.110 -83.750 ;
        RECT 69.040 -83.600 69.290 -83.490 ;
        RECT 70.790 -83.600 71.110 -83.510 ;
        RECT 69.040 -83.610 71.110 -83.600 ;
        RECT 72.580 -83.610 72.830 -83.520 ;
        RECT 73.640 -83.610 73.930 -83.560 ;
        RECT 69.040 -83.740 73.930 -83.610 ;
        RECT 69.040 -83.850 69.290 -83.740 ;
        RECT 70.790 -83.750 73.930 -83.740 ;
        RECT 70.790 -83.830 71.110 -83.750 ;
        RECT 72.580 -83.840 72.830 -83.750 ;
        RECT 73.640 -83.790 73.930 -83.750 ;
        RECT 80.860 -83.600 81.110 -83.490 ;
        RECT 82.610 -83.600 82.930 -83.510 ;
        RECT 80.860 -83.610 82.930 -83.600 ;
        RECT 84.400 -83.610 84.650 -83.520 ;
        RECT 85.460 -83.610 85.750 -83.560 ;
        RECT 80.860 -83.740 85.750 -83.610 ;
        RECT 80.860 -83.850 81.110 -83.740 ;
        RECT 82.610 -83.750 85.750 -83.740 ;
        RECT 82.610 -83.830 82.930 -83.750 ;
        RECT 84.400 -83.840 84.650 -83.750 ;
        RECT 85.460 -83.790 85.750 -83.750 ;
        RECT 92.700 -83.600 92.950 -83.490 ;
        RECT 94.450 -83.600 94.770 -83.510 ;
        RECT 92.700 -83.610 94.770 -83.600 ;
        RECT 96.240 -83.610 96.490 -83.520 ;
        RECT 97.300 -83.610 97.590 -83.560 ;
        RECT 92.700 -83.740 97.590 -83.610 ;
        RECT 92.700 -83.850 92.950 -83.740 ;
        RECT 94.450 -83.750 97.590 -83.740 ;
        RECT 94.450 -83.830 94.770 -83.750 ;
        RECT 96.240 -83.840 96.490 -83.750 ;
        RECT 97.300 -83.790 97.590 -83.750 ;
        RECT 104.540 -83.600 104.790 -83.490 ;
        RECT 106.290 -83.600 106.610 -83.510 ;
        RECT 104.540 -83.610 106.610 -83.600 ;
        RECT 108.080 -83.610 108.330 -83.520 ;
        RECT 109.140 -83.610 109.430 -83.560 ;
        RECT 104.540 -83.740 109.430 -83.610 ;
        RECT 104.540 -83.850 104.790 -83.740 ;
        RECT 106.290 -83.750 109.430 -83.740 ;
        RECT 106.290 -83.830 106.610 -83.750 ;
        RECT 108.080 -83.840 108.330 -83.750 ;
        RECT 109.140 -83.790 109.430 -83.750 ;
        RECT 116.410 -83.600 116.660 -83.490 ;
        RECT 118.160 -83.600 118.480 -83.510 ;
        RECT 116.410 -83.610 118.480 -83.600 ;
        RECT 119.950 -83.610 120.200 -83.520 ;
        RECT 121.010 -83.610 121.300 -83.560 ;
        RECT 116.410 -83.740 121.300 -83.610 ;
        RECT 116.410 -83.850 116.660 -83.740 ;
        RECT 118.160 -83.750 121.300 -83.740 ;
        RECT 118.160 -83.830 118.480 -83.750 ;
        RECT 119.950 -83.840 120.200 -83.750 ;
        RECT 121.010 -83.790 121.300 -83.750 ;
        RECT 128.280 -83.600 128.530 -83.490 ;
        RECT 130.030 -83.600 130.350 -83.510 ;
        RECT 128.280 -83.610 130.350 -83.600 ;
        RECT 131.820 -83.610 132.070 -83.520 ;
        RECT 132.880 -83.610 133.170 -83.560 ;
        RECT 128.280 -83.740 133.170 -83.610 ;
        RECT 128.280 -83.850 128.530 -83.740 ;
        RECT 130.030 -83.750 133.170 -83.740 ;
        RECT 130.030 -83.830 130.350 -83.750 ;
        RECT 131.820 -83.840 132.070 -83.750 ;
        RECT 132.880 -83.790 133.170 -83.750 ;
        RECT 137.290 -83.600 137.540 -83.490 ;
        RECT 139.040 -83.600 139.360 -83.510 ;
        RECT 137.290 -83.610 139.360 -83.600 ;
        RECT 140.830 -83.610 141.080 -83.520 ;
        RECT 141.890 -83.610 142.180 -83.560 ;
        RECT 137.290 -83.740 142.180 -83.610 ;
        RECT 137.290 -83.850 137.540 -83.740 ;
        RECT 139.040 -83.750 142.180 -83.740 ;
        RECT 139.040 -83.830 139.360 -83.750 ;
        RECT 140.830 -83.840 141.080 -83.750 ;
        RECT 141.890 -83.790 142.180 -83.750 ;
        RECT -39.910 -85.960 -39.590 -85.900 ;
        RECT -37.240 -85.950 -37.010 -85.920 ;
        RECT -33.190 -85.950 -32.960 -85.920 ;
        RECT -25.740 -85.950 -25.510 -85.920 ;
        RECT -21.690 -85.950 -21.460 -85.920 ;
        RECT -13.920 -85.950 -13.690 -85.920 ;
        RECT -9.870 -85.950 -9.640 -85.920 ;
        RECT -2.110 -85.950 -1.880 -85.920 ;
        RECT 1.940 -85.950 2.170 -85.920 ;
        RECT 9.700 -85.950 9.930 -85.920 ;
        RECT 13.750 -85.950 13.980 -85.920 ;
        RECT 21.520 -85.950 21.750 -85.920 ;
        RECT 25.570 -85.950 25.800 -85.920 ;
        RECT 33.340 -85.950 33.570 -85.920 ;
        RECT 37.390 -85.950 37.620 -85.920 ;
        RECT 45.160 -85.950 45.390 -85.920 ;
        RECT 49.210 -85.950 49.440 -85.920 ;
        RECT 56.980 -85.950 57.210 -85.920 ;
        RECT 61.030 -85.950 61.260 -85.920 ;
        RECT 68.800 -85.950 69.030 -85.920 ;
        RECT 72.850 -85.950 73.080 -85.920 ;
        RECT 80.620 -85.950 80.850 -85.920 ;
        RECT 84.670 -85.950 84.900 -85.920 ;
        RECT 92.460 -85.950 92.690 -85.920 ;
        RECT 96.510 -85.950 96.740 -85.920 ;
        RECT 104.300 -85.950 104.530 -85.920 ;
        RECT 108.350 -85.950 108.580 -85.920 ;
        RECT 116.170 -85.950 116.400 -85.920 ;
        RECT 120.220 -85.950 120.450 -85.920 ;
        RECT 128.040 -85.950 128.270 -85.920 ;
        RECT 132.090 -85.950 132.320 -85.920 ;
        RECT 137.050 -85.950 137.280 -85.920 ;
        RECT 141.100 -85.950 141.330 -85.920 ;
        RECT -37.290 -85.960 -36.960 -85.950 ;
        RECT -33.240 -85.960 -32.910 -85.950 ;
        RECT -25.790 -85.960 -25.460 -85.950 ;
        RECT -21.740 -85.960 -21.410 -85.950 ;
        RECT -13.970 -85.960 -13.640 -85.950 ;
        RECT -9.920 -85.960 -9.590 -85.950 ;
        RECT -2.160 -85.960 -1.830 -85.950 ;
        RECT 1.890 -85.960 2.220 -85.950 ;
        RECT 9.650 -85.960 9.980 -85.950 ;
        RECT 13.700 -85.960 14.030 -85.950 ;
        RECT 21.470 -85.960 21.800 -85.950 ;
        RECT 25.520 -85.960 25.850 -85.950 ;
        RECT 33.290 -85.960 33.620 -85.950 ;
        RECT 37.340 -85.960 37.670 -85.950 ;
        RECT 45.110 -85.960 45.440 -85.950 ;
        RECT 49.160 -85.960 49.490 -85.950 ;
        RECT 56.930 -85.960 57.260 -85.950 ;
        RECT 60.980 -85.960 61.310 -85.950 ;
        RECT 68.750 -85.960 69.080 -85.950 ;
        RECT 72.800 -85.960 73.130 -85.950 ;
        RECT 80.570 -85.960 80.900 -85.950 ;
        RECT 84.620 -85.960 84.950 -85.950 ;
        RECT 92.410 -85.960 92.740 -85.950 ;
        RECT 96.460 -85.960 96.790 -85.950 ;
        RECT 104.250 -85.960 104.580 -85.950 ;
        RECT 108.300 -85.960 108.630 -85.950 ;
        RECT 116.120 -85.960 116.450 -85.950 ;
        RECT 120.170 -85.960 120.500 -85.950 ;
        RECT 127.990 -85.960 128.320 -85.950 ;
        RECT 132.040 -85.960 132.370 -85.950 ;
        RECT 137.000 -85.960 137.330 -85.950 ;
        RECT 141.050 -85.960 141.380 -85.950 ;
        RECT -39.910 -86.100 142.470 -85.960 ;
        RECT -39.910 -86.160 -39.590 -86.100 ;
        RECT -37.290 -86.120 -36.960 -86.100 ;
        RECT -33.240 -86.120 -32.910 -86.100 ;
        RECT -25.790 -86.120 -25.460 -86.100 ;
        RECT -21.740 -86.120 -21.410 -86.100 ;
        RECT -13.970 -86.120 -13.640 -86.100 ;
        RECT -9.920 -86.120 -9.590 -86.100 ;
        RECT -2.160 -86.120 -1.830 -86.100 ;
        RECT 1.890 -86.120 2.220 -86.100 ;
        RECT 9.650 -86.120 9.980 -86.100 ;
        RECT 13.700 -86.120 14.030 -86.100 ;
        RECT 21.470 -86.120 21.800 -86.100 ;
        RECT 25.520 -86.120 25.850 -86.100 ;
        RECT 33.290 -86.120 33.620 -86.100 ;
        RECT 37.340 -86.120 37.670 -86.100 ;
        RECT 45.110 -86.120 45.440 -86.100 ;
        RECT 49.160 -86.120 49.490 -86.100 ;
        RECT 56.930 -86.120 57.260 -86.100 ;
        RECT 60.980 -86.120 61.310 -86.100 ;
        RECT 68.750 -86.120 69.080 -86.100 ;
        RECT 72.800 -86.120 73.130 -86.100 ;
        RECT 80.570 -86.120 80.900 -86.100 ;
        RECT 84.620 -86.120 84.950 -86.100 ;
        RECT 92.410 -86.120 92.740 -86.100 ;
        RECT 96.460 -86.120 96.790 -86.100 ;
        RECT 104.250 -86.120 104.580 -86.100 ;
        RECT 108.300 -86.120 108.630 -86.100 ;
        RECT 116.120 -86.120 116.450 -86.100 ;
        RECT 120.170 -86.120 120.500 -86.100 ;
        RECT 127.990 -86.120 128.320 -86.100 ;
        RECT 132.040 -86.120 132.370 -86.100 ;
        RECT 137.000 -86.120 137.330 -86.100 ;
        RECT 141.050 -86.120 141.380 -86.100 ;
        RECT -37.240 -86.150 -37.010 -86.120 ;
        RECT -33.190 -86.150 -32.960 -86.120 ;
        RECT -25.740 -86.150 -25.510 -86.120 ;
        RECT -21.690 -86.150 -21.460 -86.120 ;
        RECT -13.920 -86.150 -13.690 -86.120 ;
        RECT -9.870 -86.150 -9.640 -86.120 ;
        RECT -2.110 -86.150 -1.880 -86.120 ;
        RECT 1.940 -86.150 2.170 -86.120 ;
        RECT 9.700 -86.150 9.930 -86.120 ;
        RECT 13.750 -86.150 13.980 -86.120 ;
        RECT 21.520 -86.150 21.750 -86.120 ;
        RECT 25.570 -86.150 25.800 -86.120 ;
        RECT 33.340 -86.150 33.570 -86.120 ;
        RECT 37.390 -86.150 37.620 -86.120 ;
        RECT 45.160 -86.150 45.390 -86.120 ;
        RECT 49.210 -86.150 49.440 -86.120 ;
        RECT 56.980 -86.150 57.210 -86.120 ;
        RECT 61.030 -86.150 61.260 -86.120 ;
        RECT 68.800 -86.150 69.030 -86.120 ;
        RECT 72.850 -86.150 73.080 -86.120 ;
        RECT 80.620 -86.150 80.850 -86.120 ;
        RECT 84.670 -86.150 84.900 -86.120 ;
        RECT 92.460 -86.150 92.690 -86.120 ;
        RECT 96.510 -86.150 96.740 -86.120 ;
        RECT 104.300 -86.150 104.530 -86.120 ;
        RECT 108.350 -86.150 108.580 -86.120 ;
        RECT 116.170 -86.150 116.400 -86.120 ;
        RECT 120.220 -86.150 120.450 -86.120 ;
        RECT 128.040 -86.150 128.270 -86.120 ;
        RECT 132.090 -86.150 132.320 -86.120 ;
        RECT 137.050 -86.150 137.280 -86.120 ;
        RECT 141.100 -86.150 141.330 -86.120 ;
      LAYER via ;
        RECT 4.010 49.400 4.310 49.690 ;
        RECT 5.260 49.430 5.520 49.690 ;
        RECT 6.430 49.420 6.690 49.680 ;
        RECT 9.760 49.400 10.060 49.690 ;
        RECT 11.010 49.430 11.270 49.690 ;
        RECT 12.180 49.420 12.440 49.680 ;
        RECT 15.510 49.400 15.810 49.690 ;
        RECT 16.760 49.430 17.020 49.690 ;
        RECT 17.930 49.420 18.190 49.680 ;
        RECT 21.260 49.400 21.560 49.690 ;
        RECT 22.510 49.430 22.770 49.690 ;
        RECT 23.680 49.420 23.940 49.680 ;
        RECT 27.010 49.400 27.310 49.690 ;
        RECT 28.260 49.430 28.520 49.690 ;
        RECT 29.430 49.420 29.690 49.680 ;
        RECT 32.760 49.400 33.060 49.690 ;
        RECT 34.010 49.430 34.270 49.690 ;
        RECT 35.180 49.420 35.440 49.680 ;
        RECT 38.510 49.400 38.810 49.690 ;
        RECT 39.760 49.430 40.020 49.690 ;
        RECT 40.930 49.420 41.190 49.680 ;
        RECT 44.260 49.400 44.560 49.690 ;
        RECT 45.510 49.430 45.770 49.690 ;
        RECT 46.680 49.420 46.940 49.680 ;
        RECT 50.010 49.400 50.310 49.690 ;
        RECT 51.260 49.430 51.520 49.690 ;
        RECT 52.430 49.420 52.690 49.680 ;
        RECT 55.760 49.400 56.060 49.690 ;
        RECT 57.010 49.430 57.270 49.690 ;
        RECT 58.180 49.420 58.440 49.680 ;
        RECT 61.510 49.400 61.810 49.690 ;
        RECT 62.760 49.430 63.020 49.690 ;
        RECT 63.930 49.420 64.190 49.680 ;
        RECT 67.260 49.400 67.560 49.690 ;
        RECT 68.510 49.430 68.770 49.690 ;
        RECT 69.680 49.420 69.940 49.680 ;
        RECT 73.010 49.400 73.310 49.690 ;
        RECT 74.260 49.430 74.520 49.690 ;
        RECT 75.430 49.420 75.690 49.680 ;
        RECT 78.760 49.400 79.060 49.690 ;
        RECT 80.010 49.430 80.270 49.690 ;
        RECT 81.180 49.420 81.440 49.680 ;
        RECT 84.510 49.400 84.810 49.690 ;
        RECT 85.760 49.430 86.020 49.690 ;
        RECT 86.930 49.420 87.190 49.680 ;
        RECT 90.260 49.400 90.560 49.690 ;
        RECT 91.510 49.430 91.770 49.690 ;
        RECT 92.680 49.420 92.940 49.680 ;
        RECT 1.290 48.380 1.550 48.640 ;
        RECT 2.990 48.010 3.250 48.270 ;
        RECT 3.900 48.010 4.160 48.270 ;
        RECT 5.540 47.920 5.800 48.180 ;
        RECT 8.740 48.010 9.000 48.270 ;
        RECT 9.650 48.010 9.910 48.270 ;
        RECT 11.290 47.920 11.550 48.180 ;
        RECT 14.490 48.010 14.750 48.270 ;
        RECT 15.400 48.010 15.660 48.270 ;
        RECT 17.040 47.920 17.300 48.180 ;
        RECT 20.240 48.010 20.500 48.270 ;
        RECT 21.150 48.010 21.410 48.270 ;
        RECT 22.790 47.920 23.050 48.180 ;
        RECT 25.990 48.010 26.250 48.270 ;
        RECT 26.900 48.010 27.160 48.270 ;
        RECT 28.540 47.920 28.800 48.180 ;
        RECT 31.740 48.010 32.000 48.270 ;
        RECT 32.650 48.010 32.910 48.270 ;
        RECT 34.290 47.920 34.550 48.180 ;
        RECT 37.490 48.010 37.750 48.270 ;
        RECT 38.400 48.010 38.660 48.270 ;
        RECT 40.040 47.920 40.300 48.180 ;
        RECT 43.240 48.010 43.500 48.270 ;
        RECT 44.150 48.010 44.410 48.270 ;
        RECT 45.790 47.920 46.050 48.180 ;
        RECT 48.990 48.010 49.250 48.270 ;
        RECT 49.900 48.010 50.160 48.270 ;
        RECT 51.540 47.920 51.800 48.180 ;
        RECT 54.740 48.010 55.000 48.270 ;
        RECT 55.650 48.010 55.910 48.270 ;
        RECT 57.290 47.920 57.550 48.180 ;
        RECT 60.490 48.010 60.750 48.270 ;
        RECT 61.400 48.010 61.660 48.270 ;
        RECT 63.040 47.920 63.300 48.180 ;
        RECT 66.240 48.010 66.500 48.270 ;
        RECT 67.150 48.010 67.410 48.270 ;
        RECT 68.790 47.920 69.050 48.180 ;
        RECT 71.990 48.010 72.250 48.270 ;
        RECT 72.900 48.010 73.160 48.270 ;
        RECT 74.540 47.920 74.800 48.180 ;
        RECT 77.740 48.010 78.000 48.270 ;
        RECT 78.650 48.010 78.910 48.270 ;
        RECT 80.290 47.920 80.550 48.180 ;
        RECT 83.490 48.010 83.750 48.270 ;
        RECT 84.400 48.010 84.660 48.270 ;
        RECT 86.040 47.920 86.300 48.180 ;
        RECT 89.240 48.010 89.500 48.270 ;
        RECT 90.150 48.010 90.410 48.270 ;
        RECT 91.790 47.920 92.050 48.180 ;
        RECT 1.280 47.550 1.540 47.810 ;
        RECT 1.300 46.690 1.560 46.950 ;
        RECT 1.280 45.970 1.540 46.230 ;
        RECT 4.960 46.330 5.220 46.590 ;
        RECT 6.600 46.330 6.860 46.590 ;
        RECT 7.510 46.330 7.770 46.590 ;
        RECT 10.710 46.330 10.970 46.590 ;
        RECT 12.350 46.330 12.610 46.590 ;
        RECT 13.260 46.330 13.520 46.590 ;
        RECT 16.460 46.330 16.720 46.590 ;
        RECT 18.100 46.330 18.360 46.590 ;
        RECT 19.010 46.330 19.270 46.590 ;
        RECT 22.210 46.330 22.470 46.590 ;
        RECT 23.850 46.330 24.110 46.590 ;
        RECT 24.760 46.330 25.020 46.590 ;
        RECT 27.960 46.330 28.220 46.590 ;
        RECT 29.600 46.330 29.860 46.590 ;
        RECT 30.510 46.330 30.770 46.590 ;
        RECT 33.710 46.330 33.970 46.590 ;
        RECT 35.350 46.330 35.610 46.590 ;
        RECT 36.260 46.330 36.520 46.590 ;
        RECT 39.460 46.330 39.720 46.590 ;
        RECT 41.100 46.330 41.360 46.590 ;
        RECT 42.010 46.330 42.270 46.590 ;
        RECT 45.210 46.330 45.470 46.590 ;
        RECT 46.850 46.330 47.110 46.590 ;
        RECT 47.760 46.330 48.020 46.590 ;
        RECT 50.960 46.330 51.220 46.590 ;
        RECT 52.600 46.330 52.860 46.590 ;
        RECT 53.510 46.330 53.770 46.590 ;
        RECT 56.710 46.330 56.970 46.590 ;
        RECT 58.350 46.330 58.610 46.590 ;
        RECT 59.260 46.330 59.520 46.590 ;
        RECT 62.460 46.330 62.720 46.590 ;
        RECT 64.100 46.330 64.360 46.590 ;
        RECT 65.010 46.330 65.270 46.590 ;
        RECT 68.210 46.330 68.470 46.590 ;
        RECT 69.850 46.330 70.110 46.590 ;
        RECT 70.760 46.330 71.020 46.590 ;
        RECT 73.960 46.330 74.220 46.590 ;
        RECT 75.600 46.330 75.860 46.590 ;
        RECT 76.510 46.330 76.770 46.590 ;
        RECT 79.710 46.330 79.970 46.590 ;
        RECT 81.350 46.330 81.610 46.590 ;
        RECT 82.260 46.330 82.520 46.590 ;
        RECT 85.460 46.330 85.720 46.590 ;
        RECT 87.100 46.330 87.360 46.590 ;
        RECT 88.010 46.330 88.270 46.590 ;
        RECT 91.210 46.330 91.470 46.590 ;
        RECT 92.850 46.330 93.110 46.590 ;
        RECT 93.760 46.330 94.020 46.590 ;
        RECT 2.990 45.600 3.250 45.860 ;
        RECT 3.900 45.600 4.160 45.860 ;
        RECT 5.540 45.510 5.800 45.770 ;
        RECT 8.740 45.600 9.000 45.860 ;
        RECT 9.650 45.600 9.910 45.860 ;
        RECT 11.290 45.510 11.550 45.770 ;
        RECT 14.490 45.600 14.750 45.860 ;
        RECT 15.400 45.600 15.660 45.860 ;
        RECT 17.040 45.510 17.300 45.770 ;
        RECT 20.240 45.600 20.500 45.860 ;
        RECT 21.150 45.600 21.410 45.860 ;
        RECT 22.790 45.510 23.050 45.770 ;
        RECT 25.990 45.600 26.250 45.860 ;
        RECT 26.900 45.600 27.160 45.860 ;
        RECT 28.540 45.510 28.800 45.770 ;
        RECT 31.740 45.600 32.000 45.860 ;
        RECT 32.650 45.600 32.910 45.860 ;
        RECT 34.290 45.510 34.550 45.770 ;
        RECT 37.490 45.600 37.750 45.860 ;
        RECT 38.400 45.600 38.660 45.860 ;
        RECT 40.040 45.510 40.300 45.770 ;
        RECT 43.240 45.600 43.500 45.860 ;
        RECT 44.150 45.600 44.410 45.860 ;
        RECT 45.790 45.510 46.050 45.770 ;
        RECT 48.990 45.600 49.250 45.860 ;
        RECT 49.900 45.600 50.160 45.860 ;
        RECT 51.540 45.510 51.800 45.770 ;
        RECT 54.740 45.600 55.000 45.860 ;
        RECT 55.650 45.600 55.910 45.860 ;
        RECT 57.290 45.510 57.550 45.770 ;
        RECT 60.490 45.600 60.750 45.860 ;
        RECT 61.400 45.600 61.660 45.860 ;
        RECT 63.040 45.510 63.300 45.770 ;
        RECT 66.240 45.600 66.500 45.860 ;
        RECT 67.150 45.600 67.410 45.860 ;
        RECT 68.790 45.510 69.050 45.770 ;
        RECT 71.990 45.600 72.250 45.860 ;
        RECT 72.900 45.600 73.160 45.860 ;
        RECT 74.540 45.510 74.800 45.770 ;
        RECT 77.740 45.600 78.000 45.860 ;
        RECT 78.650 45.600 78.910 45.860 ;
        RECT 80.290 45.510 80.550 45.770 ;
        RECT 83.490 45.600 83.750 45.860 ;
        RECT 84.400 45.600 84.660 45.860 ;
        RECT 86.040 45.510 86.300 45.770 ;
        RECT 89.240 45.600 89.500 45.860 ;
        RECT 90.150 45.600 90.410 45.860 ;
        RECT 91.790 45.510 92.050 45.770 ;
        RECT 1.290 45.120 1.550 45.380 ;
        RECT 1.290 44.320 1.550 44.580 ;
        RECT 1.280 43.560 1.540 43.820 ;
        RECT 4.960 43.920 5.220 44.180 ;
        RECT 6.600 43.920 6.860 44.180 ;
        RECT 7.510 43.920 7.770 44.180 ;
        RECT 10.710 43.920 10.970 44.180 ;
        RECT 12.350 43.920 12.610 44.180 ;
        RECT 13.260 43.920 13.520 44.180 ;
        RECT 16.460 43.920 16.720 44.180 ;
        RECT 18.100 43.920 18.360 44.180 ;
        RECT 19.010 43.920 19.270 44.180 ;
        RECT 22.210 43.920 22.470 44.180 ;
        RECT 23.850 43.920 24.110 44.180 ;
        RECT 24.760 43.920 25.020 44.180 ;
        RECT 27.960 43.920 28.220 44.180 ;
        RECT 29.600 43.920 29.860 44.180 ;
        RECT 30.510 43.920 30.770 44.180 ;
        RECT 33.710 43.920 33.970 44.180 ;
        RECT 35.350 43.920 35.610 44.180 ;
        RECT 36.260 43.920 36.520 44.180 ;
        RECT 39.460 43.920 39.720 44.180 ;
        RECT 41.100 43.920 41.360 44.180 ;
        RECT 42.010 43.920 42.270 44.180 ;
        RECT 45.210 43.920 45.470 44.180 ;
        RECT 46.850 43.920 47.110 44.180 ;
        RECT 47.760 43.920 48.020 44.180 ;
        RECT 50.960 43.920 51.220 44.180 ;
        RECT 52.600 43.920 52.860 44.180 ;
        RECT 53.510 43.920 53.770 44.180 ;
        RECT 56.710 43.920 56.970 44.180 ;
        RECT 58.350 43.920 58.610 44.180 ;
        RECT 59.260 43.920 59.520 44.180 ;
        RECT 62.460 43.920 62.720 44.180 ;
        RECT 64.100 43.920 64.360 44.180 ;
        RECT 65.010 43.920 65.270 44.180 ;
        RECT 68.210 43.920 68.470 44.180 ;
        RECT 69.850 43.920 70.110 44.180 ;
        RECT 70.760 43.920 71.020 44.180 ;
        RECT 73.960 43.920 74.220 44.180 ;
        RECT 75.600 43.920 75.860 44.180 ;
        RECT 76.510 43.920 76.770 44.180 ;
        RECT 79.710 43.920 79.970 44.180 ;
        RECT 81.350 43.920 81.610 44.180 ;
        RECT 82.260 43.920 82.520 44.180 ;
        RECT 85.460 43.920 85.720 44.180 ;
        RECT 87.100 43.920 87.360 44.180 ;
        RECT 88.010 43.920 88.270 44.180 ;
        RECT 91.210 43.920 91.470 44.180 ;
        RECT 92.850 43.920 93.110 44.180 ;
        RECT 93.760 43.920 94.020 44.180 ;
        RECT 2.990 42.630 3.250 42.890 ;
        RECT 3.900 42.630 4.160 42.890 ;
        RECT 5.540 42.540 5.800 42.800 ;
        RECT 8.740 42.630 9.000 42.890 ;
        RECT 9.650 42.630 9.910 42.890 ;
        RECT 11.290 42.540 11.550 42.800 ;
        RECT 14.490 42.630 14.750 42.890 ;
        RECT 15.400 42.630 15.660 42.890 ;
        RECT 17.040 42.540 17.300 42.800 ;
        RECT 20.240 42.630 20.500 42.890 ;
        RECT 21.150 42.630 21.410 42.890 ;
        RECT 22.790 42.540 23.050 42.800 ;
        RECT 25.990 42.630 26.250 42.890 ;
        RECT 26.900 42.630 27.160 42.890 ;
        RECT 28.540 42.540 28.800 42.800 ;
        RECT 31.740 42.630 32.000 42.890 ;
        RECT 32.650 42.630 32.910 42.890 ;
        RECT 34.290 42.540 34.550 42.800 ;
        RECT 37.490 42.630 37.750 42.890 ;
        RECT 38.400 42.630 38.660 42.890 ;
        RECT 40.040 42.540 40.300 42.800 ;
        RECT 43.240 42.630 43.500 42.890 ;
        RECT 44.150 42.630 44.410 42.890 ;
        RECT 45.790 42.540 46.050 42.800 ;
        RECT 48.990 42.630 49.250 42.890 ;
        RECT 49.900 42.630 50.160 42.890 ;
        RECT 51.540 42.540 51.800 42.800 ;
        RECT 54.740 42.630 55.000 42.890 ;
        RECT 55.650 42.630 55.910 42.890 ;
        RECT 57.290 42.540 57.550 42.800 ;
        RECT 60.490 42.630 60.750 42.890 ;
        RECT 61.400 42.630 61.660 42.890 ;
        RECT 63.040 42.540 63.300 42.800 ;
        RECT 66.240 42.630 66.500 42.890 ;
        RECT 67.150 42.630 67.410 42.890 ;
        RECT 68.790 42.540 69.050 42.800 ;
        RECT 71.990 42.630 72.250 42.890 ;
        RECT 72.900 42.630 73.160 42.890 ;
        RECT 74.540 42.540 74.800 42.800 ;
        RECT 77.740 42.630 78.000 42.890 ;
        RECT 78.650 42.630 78.910 42.890 ;
        RECT 80.290 42.540 80.550 42.800 ;
        RECT 83.490 42.630 83.750 42.890 ;
        RECT 84.400 42.630 84.660 42.890 ;
        RECT 86.040 42.540 86.300 42.800 ;
        RECT 89.240 42.630 89.500 42.890 ;
        RECT 90.150 42.630 90.410 42.890 ;
        RECT 91.790 42.540 92.050 42.800 ;
        RECT 1.300 42.190 1.560 42.450 ;
        RECT 1.300 41.330 1.560 41.590 ;
        RECT 1.280 40.590 1.540 40.850 ;
        RECT 4.960 40.950 5.220 41.210 ;
        RECT 6.600 40.950 6.860 41.210 ;
        RECT 7.510 40.950 7.770 41.210 ;
        RECT 10.710 40.950 10.970 41.210 ;
        RECT 12.350 40.950 12.610 41.210 ;
        RECT 13.260 40.950 13.520 41.210 ;
        RECT 16.460 40.950 16.720 41.210 ;
        RECT 18.100 40.950 18.360 41.210 ;
        RECT 19.010 40.950 19.270 41.210 ;
        RECT 22.210 40.950 22.470 41.210 ;
        RECT 23.850 40.950 24.110 41.210 ;
        RECT 24.760 40.950 25.020 41.210 ;
        RECT 27.960 40.950 28.220 41.210 ;
        RECT 29.600 40.950 29.860 41.210 ;
        RECT 30.510 40.950 30.770 41.210 ;
        RECT 33.710 40.950 33.970 41.210 ;
        RECT 35.350 40.950 35.610 41.210 ;
        RECT 36.260 40.950 36.520 41.210 ;
        RECT 39.460 40.950 39.720 41.210 ;
        RECT 41.100 40.950 41.360 41.210 ;
        RECT 42.010 40.950 42.270 41.210 ;
        RECT 45.210 40.950 45.470 41.210 ;
        RECT 46.850 40.950 47.110 41.210 ;
        RECT 47.760 40.950 48.020 41.210 ;
        RECT 50.960 40.950 51.220 41.210 ;
        RECT 52.600 40.950 52.860 41.210 ;
        RECT 53.510 40.950 53.770 41.210 ;
        RECT 56.710 40.950 56.970 41.210 ;
        RECT 58.350 40.950 58.610 41.210 ;
        RECT 59.260 40.950 59.520 41.210 ;
        RECT 62.460 40.950 62.720 41.210 ;
        RECT 64.100 40.950 64.360 41.210 ;
        RECT 65.010 40.950 65.270 41.210 ;
        RECT 68.210 40.950 68.470 41.210 ;
        RECT 69.850 40.950 70.110 41.210 ;
        RECT 70.760 40.950 71.020 41.210 ;
        RECT 73.960 40.950 74.220 41.210 ;
        RECT 75.600 40.950 75.860 41.210 ;
        RECT 76.510 40.950 76.770 41.210 ;
        RECT 79.710 40.950 79.970 41.210 ;
        RECT 81.350 40.950 81.610 41.210 ;
        RECT 82.260 40.950 82.520 41.210 ;
        RECT 85.460 40.950 85.720 41.210 ;
        RECT 87.100 40.950 87.360 41.210 ;
        RECT 88.010 40.950 88.270 41.210 ;
        RECT 91.210 40.950 91.470 41.210 ;
        RECT 92.850 40.950 93.110 41.210 ;
        RECT 93.760 40.950 94.020 41.210 ;
        RECT 2.990 40.220 3.250 40.480 ;
        RECT 3.900 40.220 4.160 40.480 ;
        RECT 5.540 40.130 5.800 40.390 ;
        RECT 8.740 40.220 9.000 40.480 ;
        RECT 9.650 40.220 9.910 40.480 ;
        RECT 11.290 40.130 11.550 40.390 ;
        RECT 14.490 40.220 14.750 40.480 ;
        RECT 15.400 40.220 15.660 40.480 ;
        RECT 17.040 40.130 17.300 40.390 ;
        RECT 20.240 40.220 20.500 40.480 ;
        RECT 21.150 40.220 21.410 40.480 ;
        RECT 22.790 40.130 23.050 40.390 ;
        RECT 25.990 40.220 26.250 40.480 ;
        RECT 26.900 40.220 27.160 40.480 ;
        RECT 28.540 40.130 28.800 40.390 ;
        RECT 31.740 40.220 32.000 40.480 ;
        RECT 32.650 40.220 32.910 40.480 ;
        RECT 34.290 40.130 34.550 40.390 ;
        RECT 37.490 40.220 37.750 40.480 ;
        RECT 38.400 40.220 38.660 40.480 ;
        RECT 40.040 40.130 40.300 40.390 ;
        RECT 43.240 40.220 43.500 40.480 ;
        RECT 44.150 40.220 44.410 40.480 ;
        RECT 45.790 40.130 46.050 40.390 ;
        RECT 48.990 40.220 49.250 40.480 ;
        RECT 49.900 40.220 50.160 40.480 ;
        RECT 51.540 40.130 51.800 40.390 ;
        RECT 54.740 40.220 55.000 40.480 ;
        RECT 55.650 40.220 55.910 40.480 ;
        RECT 57.290 40.130 57.550 40.390 ;
        RECT 60.490 40.220 60.750 40.480 ;
        RECT 61.400 40.220 61.660 40.480 ;
        RECT 63.040 40.130 63.300 40.390 ;
        RECT 66.240 40.220 66.500 40.480 ;
        RECT 67.150 40.220 67.410 40.480 ;
        RECT 68.790 40.130 69.050 40.390 ;
        RECT 71.990 40.220 72.250 40.480 ;
        RECT 72.900 40.220 73.160 40.480 ;
        RECT 74.540 40.130 74.800 40.390 ;
        RECT 77.740 40.220 78.000 40.480 ;
        RECT 78.650 40.220 78.910 40.480 ;
        RECT 80.290 40.130 80.550 40.390 ;
        RECT 83.490 40.220 83.750 40.480 ;
        RECT 84.400 40.220 84.660 40.480 ;
        RECT 86.040 40.130 86.300 40.390 ;
        RECT 89.240 40.220 89.500 40.480 ;
        RECT 90.150 40.220 90.410 40.480 ;
        RECT 91.790 40.130 92.050 40.390 ;
        RECT 1.300 39.760 1.560 40.020 ;
        RECT 1.300 38.920 1.560 39.180 ;
        RECT 1.290 38.180 1.550 38.440 ;
        RECT 4.960 38.540 5.220 38.800 ;
        RECT 6.600 38.540 6.860 38.800 ;
        RECT 7.510 38.540 7.770 38.800 ;
        RECT 10.710 38.540 10.970 38.800 ;
        RECT 12.350 38.540 12.610 38.800 ;
        RECT 13.260 38.540 13.520 38.800 ;
        RECT 16.460 38.540 16.720 38.800 ;
        RECT 18.100 38.540 18.360 38.800 ;
        RECT 19.010 38.540 19.270 38.800 ;
        RECT 22.210 38.540 22.470 38.800 ;
        RECT 23.850 38.540 24.110 38.800 ;
        RECT 24.760 38.540 25.020 38.800 ;
        RECT 27.960 38.540 28.220 38.800 ;
        RECT 29.600 38.540 29.860 38.800 ;
        RECT 30.510 38.540 30.770 38.800 ;
        RECT 33.710 38.540 33.970 38.800 ;
        RECT 35.350 38.540 35.610 38.800 ;
        RECT 36.260 38.540 36.520 38.800 ;
        RECT 39.460 38.540 39.720 38.800 ;
        RECT 41.100 38.540 41.360 38.800 ;
        RECT 42.010 38.540 42.270 38.800 ;
        RECT 45.210 38.540 45.470 38.800 ;
        RECT 46.850 38.540 47.110 38.800 ;
        RECT 47.760 38.540 48.020 38.800 ;
        RECT 50.960 38.540 51.220 38.800 ;
        RECT 52.600 38.540 52.860 38.800 ;
        RECT 53.510 38.540 53.770 38.800 ;
        RECT 56.710 38.540 56.970 38.800 ;
        RECT 58.350 38.540 58.610 38.800 ;
        RECT 59.260 38.540 59.520 38.800 ;
        RECT 62.460 38.540 62.720 38.800 ;
        RECT 64.100 38.540 64.360 38.800 ;
        RECT 65.010 38.540 65.270 38.800 ;
        RECT 68.210 38.540 68.470 38.800 ;
        RECT 69.850 38.540 70.110 38.800 ;
        RECT 70.760 38.540 71.020 38.800 ;
        RECT 73.960 38.540 74.220 38.800 ;
        RECT 75.600 38.540 75.860 38.800 ;
        RECT 76.510 38.540 76.770 38.800 ;
        RECT 79.710 38.540 79.970 38.800 ;
        RECT 81.350 38.540 81.610 38.800 ;
        RECT 82.260 38.540 82.520 38.800 ;
        RECT 85.460 38.540 85.720 38.800 ;
        RECT 87.100 38.540 87.360 38.800 ;
        RECT 88.010 38.540 88.270 38.800 ;
        RECT 91.210 38.540 91.470 38.800 ;
        RECT 92.850 38.540 93.110 38.800 ;
        RECT 93.760 38.540 94.020 38.800 ;
        RECT 2.990 37.810 3.250 38.070 ;
        RECT 3.900 37.810 4.160 38.070 ;
        RECT 5.540 37.720 5.800 37.980 ;
        RECT 8.740 37.810 9.000 38.070 ;
        RECT 9.650 37.810 9.910 38.070 ;
        RECT 11.290 37.720 11.550 37.980 ;
        RECT 14.490 37.810 14.750 38.070 ;
        RECT 15.400 37.810 15.660 38.070 ;
        RECT 17.040 37.720 17.300 37.980 ;
        RECT 20.240 37.810 20.500 38.070 ;
        RECT 21.150 37.810 21.410 38.070 ;
        RECT 22.790 37.720 23.050 37.980 ;
        RECT 25.990 37.810 26.250 38.070 ;
        RECT 26.900 37.810 27.160 38.070 ;
        RECT 28.540 37.720 28.800 37.980 ;
        RECT 31.740 37.810 32.000 38.070 ;
        RECT 32.650 37.810 32.910 38.070 ;
        RECT 34.290 37.720 34.550 37.980 ;
        RECT 37.490 37.810 37.750 38.070 ;
        RECT 38.400 37.810 38.660 38.070 ;
        RECT 40.040 37.720 40.300 37.980 ;
        RECT 43.240 37.810 43.500 38.070 ;
        RECT 44.150 37.810 44.410 38.070 ;
        RECT 45.790 37.720 46.050 37.980 ;
        RECT 48.990 37.810 49.250 38.070 ;
        RECT 49.900 37.810 50.160 38.070 ;
        RECT 51.540 37.720 51.800 37.980 ;
        RECT 54.740 37.810 55.000 38.070 ;
        RECT 55.650 37.810 55.910 38.070 ;
        RECT 57.290 37.720 57.550 37.980 ;
        RECT 60.490 37.810 60.750 38.070 ;
        RECT 61.400 37.810 61.660 38.070 ;
        RECT 63.040 37.720 63.300 37.980 ;
        RECT 66.240 37.810 66.500 38.070 ;
        RECT 67.150 37.810 67.410 38.070 ;
        RECT 68.790 37.720 69.050 37.980 ;
        RECT 71.990 37.810 72.250 38.070 ;
        RECT 72.900 37.810 73.160 38.070 ;
        RECT 74.540 37.720 74.800 37.980 ;
        RECT 77.740 37.810 78.000 38.070 ;
        RECT 78.650 37.810 78.910 38.070 ;
        RECT 80.290 37.720 80.550 37.980 ;
        RECT 83.490 37.810 83.750 38.070 ;
        RECT 84.400 37.810 84.660 38.070 ;
        RECT 86.040 37.720 86.300 37.980 ;
        RECT 89.240 37.810 89.500 38.070 ;
        RECT 90.150 37.810 90.410 38.070 ;
        RECT 91.790 37.720 92.050 37.980 ;
        RECT 1.290 35.770 1.550 36.030 ;
        RECT 4.960 36.130 5.220 36.390 ;
        RECT 6.600 36.130 6.860 36.390 ;
        RECT 7.510 36.130 7.770 36.390 ;
        RECT 10.710 36.130 10.970 36.390 ;
        RECT 12.350 36.130 12.610 36.390 ;
        RECT 13.260 36.130 13.520 36.390 ;
        RECT 16.460 36.130 16.720 36.390 ;
        RECT 18.100 36.130 18.360 36.390 ;
        RECT 19.010 36.130 19.270 36.390 ;
        RECT 22.210 36.130 22.470 36.390 ;
        RECT 23.850 36.130 24.110 36.390 ;
        RECT 24.760 36.130 25.020 36.390 ;
        RECT 27.960 36.130 28.220 36.390 ;
        RECT 29.600 36.130 29.860 36.390 ;
        RECT 30.510 36.130 30.770 36.390 ;
        RECT 33.710 36.130 33.970 36.390 ;
        RECT 35.350 36.130 35.610 36.390 ;
        RECT 36.260 36.130 36.520 36.390 ;
        RECT 39.460 36.130 39.720 36.390 ;
        RECT 41.100 36.130 41.360 36.390 ;
        RECT 42.010 36.130 42.270 36.390 ;
        RECT 45.210 36.130 45.470 36.390 ;
        RECT 46.850 36.130 47.110 36.390 ;
        RECT 47.760 36.130 48.020 36.390 ;
        RECT 50.960 36.130 51.220 36.390 ;
        RECT 52.600 36.130 52.860 36.390 ;
        RECT 53.510 36.130 53.770 36.390 ;
        RECT 56.710 36.130 56.970 36.390 ;
        RECT 58.350 36.130 58.610 36.390 ;
        RECT 59.260 36.130 59.520 36.390 ;
        RECT 62.460 36.130 62.720 36.390 ;
        RECT 64.100 36.130 64.360 36.390 ;
        RECT 65.010 36.130 65.270 36.390 ;
        RECT 68.210 36.130 68.470 36.390 ;
        RECT 69.850 36.130 70.110 36.390 ;
        RECT 70.760 36.130 71.020 36.390 ;
        RECT 73.960 36.130 74.220 36.390 ;
        RECT 75.600 36.130 75.860 36.390 ;
        RECT 76.510 36.130 76.770 36.390 ;
        RECT 79.710 36.130 79.970 36.390 ;
        RECT 81.350 36.130 81.610 36.390 ;
        RECT 82.260 36.130 82.520 36.390 ;
        RECT 85.460 36.130 85.720 36.390 ;
        RECT 87.100 36.130 87.360 36.390 ;
        RECT 88.010 36.130 88.270 36.390 ;
        RECT 91.210 36.130 91.470 36.390 ;
        RECT 92.850 36.130 93.110 36.390 ;
        RECT 93.760 36.130 94.020 36.390 ;
        RECT 2.990 35.400 3.250 35.660 ;
        RECT 3.900 35.400 4.160 35.660 ;
        RECT 5.540 35.310 5.800 35.570 ;
        RECT 8.740 35.400 9.000 35.660 ;
        RECT 9.650 35.400 9.910 35.660 ;
        RECT 11.290 35.310 11.550 35.570 ;
        RECT 14.490 35.400 14.750 35.660 ;
        RECT 15.400 35.400 15.660 35.660 ;
        RECT 17.040 35.310 17.300 35.570 ;
        RECT 20.240 35.400 20.500 35.660 ;
        RECT 21.150 35.400 21.410 35.660 ;
        RECT 22.790 35.310 23.050 35.570 ;
        RECT 25.990 35.400 26.250 35.660 ;
        RECT 26.900 35.400 27.160 35.660 ;
        RECT 28.540 35.310 28.800 35.570 ;
        RECT 31.740 35.400 32.000 35.660 ;
        RECT 32.650 35.400 32.910 35.660 ;
        RECT 34.290 35.310 34.550 35.570 ;
        RECT 37.490 35.400 37.750 35.660 ;
        RECT 38.400 35.400 38.660 35.660 ;
        RECT 40.040 35.310 40.300 35.570 ;
        RECT 43.240 35.400 43.500 35.660 ;
        RECT 44.150 35.400 44.410 35.660 ;
        RECT 45.790 35.310 46.050 35.570 ;
        RECT 48.990 35.400 49.250 35.660 ;
        RECT 49.900 35.400 50.160 35.660 ;
        RECT 51.540 35.310 51.800 35.570 ;
        RECT 54.740 35.400 55.000 35.660 ;
        RECT 55.650 35.400 55.910 35.660 ;
        RECT 57.290 35.310 57.550 35.570 ;
        RECT 60.490 35.400 60.750 35.660 ;
        RECT 61.400 35.400 61.660 35.660 ;
        RECT 63.040 35.310 63.300 35.570 ;
        RECT 66.240 35.400 66.500 35.660 ;
        RECT 67.150 35.400 67.410 35.660 ;
        RECT 68.790 35.310 69.050 35.570 ;
        RECT 71.990 35.400 72.250 35.660 ;
        RECT 72.900 35.400 73.160 35.660 ;
        RECT 74.540 35.310 74.800 35.570 ;
        RECT 77.740 35.400 78.000 35.660 ;
        RECT 78.650 35.400 78.910 35.660 ;
        RECT 80.290 35.310 80.550 35.570 ;
        RECT 83.490 35.400 83.750 35.660 ;
        RECT 84.400 35.400 84.660 35.660 ;
        RECT 86.040 35.310 86.300 35.570 ;
        RECT 89.240 35.400 89.500 35.660 ;
        RECT 90.150 35.400 90.410 35.660 ;
        RECT 91.790 35.310 92.050 35.570 ;
        RECT 1.290 33.360 1.550 33.620 ;
        RECT 4.960 33.720 5.220 33.980 ;
        RECT 6.600 33.720 6.860 33.980 ;
        RECT 7.510 33.720 7.770 33.980 ;
        RECT 10.710 33.720 10.970 33.980 ;
        RECT 12.350 33.720 12.610 33.980 ;
        RECT 13.260 33.720 13.520 33.980 ;
        RECT 16.460 33.720 16.720 33.980 ;
        RECT 18.100 33.720 18.360 33.980 ;
        RECT 19.010 33.720 19.270 33.980 ;
        RECT 22.210 33.720 22.470 33.980 ;
        RECT 23.850 33.720 24.110 33.980 ;
        RECT 24.760 33.720 25.020 33.980 ;
        RECT 27.960 33.720 28.220 33.980 ;
        RECT 29.600 33.720 29.860 33.980 ;
        RECT 30.510 33.720 30.770 33.980 ;
        RECT 33.710 33.720 33.970 33.980 ;
        RECT 35.350 33.720 35.610 33.980 ;
        RECT 36.260 33.720 36.520 33.980 ;
        RECT 39.460 33.720 39.720 33.980 ;
        RECT 41.100 33.720 41.360 33.980 ;
        RECT 42.010 33.720 42.270 33.980 ;
        RECT 45.210 33.720 45.470 33.980 ;
        RECT 46.850 33.720 47.110 33.980 ;
        RECT 47.760 33.720 48.020 33.980 ;
        RECT 50.960 33.720 51.220 33.980 ;
        RECT 52.600 33.720 52.860 33.980 ;
        RECT 53.510 33.720 53.770 33.980 ;
        RECT 56.710 33.720 56.970 33.980 ;
        RECT 58.350 33.720 58.610 33.980 ;
        RECT 59.260 33.720 59.520 33.980 ;
        RECT 62.460 33.720 62.720 33.980 ;
        RECT 64.100 33.720 64.360 33.980 ;
        RECT 65.010 33.720 65.270 33.980 ;
        RECT 68.210 33.720 68.470 33.980 ;
        RECT 69.850 33.720 70.110 33.980 ;
        RECT 70.760 33.720 71.020 33.980 ;
        RECT 73.960 33.720 74.220 33.980 ;
        RECT 75.600 33.720 75.860 33.980 ;
        RECT 76.510 33.720 76.770 33.980 ;
        RECT 79.710 33.720 79.970 33.980 ;
        RECT 81.350 33.720 81.610 33.980 ;
        RECT 82.260 33.720 82.520 33.980 ;
        RECT 85.460 33.720 85.720 33.980 ;
        RECT 87.100 33.720 87.360 33.980 ;
        RECT 88.010 33.720 88.270 33.980 ;
        RECT 91.210 33.720 91.470 33.980 ;
        RECT 92.850 33.720 93.110 33.980 ;
        RECT 93.760 33.720 94.020 33.980 ;
        RECT 2.990 32.990 3.250 33.250 ;
        RECT 3.900 32.990 4.160 33.250 ;
        RECT 5.540 32.900 5.800 33.160 ;
        RECT 8.740 32.990 9.000 33.250 ;
        RECT 9.650 32.990 9.910 33.250 ;
        RECT 11.290 32.900 11.550 33.160 ;
        RECT 14.490 32.990 14.750 33.250 ;
        RECT 15.400 32.990 15.660 33.250 ;
        RECT 17.040 32.900 17.300 33.160 ;
        RECT 20.240 32.990 20.500 33.250 ;
        RECT 21.150 32.990 21.410 33.250 ;
        RECT 22.790 32.900 23.050 33.160 ;
        RECT 25.990 32.990 26.250 33.250 ;
        RECT 26.900 32.990 27.160 33.250 ;
        RECT 28.540 32.900 28.800 33.160 ;
        RECT 31.740 32.990 32.000 33.250 ;
        RECT 32.650 32.990 32.910 33.250 ;
        RECT 34.290 32.900 34.550 33.160 ;
        RECT 37.490 32.990 37.750 33.250 ;
        RECT 38.400 32.990 38.660 33.250 ;
        RECT 40.040 32.900 40.300 33.160 ;
        RECT 43.240 32.990 43.500 33.250 ;
        RECT 44.150 32.990 44.410 33.250 ;
        RECT 45.790 32.900 46.050 33.160 ;
        RECT 48.990 32.990 49.250 33.250 ;
        RECT 49.900 32.990 50.160 33.250 ;
        RECT 51.540 32.900 51.800 33.160 ;
        RECT 54.740 32.990 55.000 33.250 ;
        RECT 55.650 32.990 55.910 33.250 ;
        RECT 57.290 32.900 57.550 33.160 ;
        RECT 60.490 32.990 60.750 33.250 ;
        RECT 61.400 32.990 61.660 33.250 ;
        RECT 63.040 32.900 63.300 33.160 ;
        RECT 66.240 32.990 66.500 33.250 ;
        RECT 67.150 32.990 67.410 33.250 ;
        RECT 68.790 32.900 69.050 33.160 ;
        RECT 71.990 32.990 72.250 33.250 ;
        RECT 72.900 32.990 73.160 33.250 ;
        RECT 74.540 32.900 74.800 33.160 ;
        RECT 77.740 32.990 78.000 33.250 ;
        RECT 78.650 32.990 78.910 33.250 ;
        RECT 80.290 32.900 80.550 33.160 ;
        RECT 83.490 32.990 83.750 33.250 ;
        RECT 84.400 32.990 84.660 33.250 ;
        RECT 86.040 32.900 86.300 33.160 ;
        RECT 89.240 32.990 89.500 33.250 ;
        RECT 90.150 32.990 90.410 33.250 ;
        RECT 91.790 32.900 92.050 33.160 ;
        RECT 1.290 30.950 1.550 31.210 ;
        RECT 4.960 31.310 5.220 31.570 ;
        RECT 6.600 31.310 6.860 31.570 ;
        RECT 7.510 31.310 7.770 31.570 ;
        RECT 10.710 31.310 10.970 31.570 ;
        RECT 12.350 31.310 12.610 31.570 ;
        RECT 13.260 31.310 13.520 31.570 ;
        RECT 16.460 31.310 16.720 31.570 ;
        RECT 18.100 31.310 18.360 31.570 ;
        RECT 19.010 31.310 19.270 31.570 ;
        RECT 22.210 31.310 22.470 31.570 ;
        RECT 23.850 31.310 24.110 31.570 ;
        RECT 24.760 31.310 25.020 31.570 ;
        RECT 27.960 31.310 28.220 31.570 ;
        RECT 29.600 31.310 29.860 31.570 ;
        RECT 30.510 31.310 30.770 31.570 ;
        RECT 33.710 31.310 33.970 31.570 ;
        RECT 35.350 31.310 35.610 31.570 ;
        RECT 36.260 31.310 36.520 31.570 ;
        RECT 39.460 31.310 39.720 31.570 ;
        RECT 41.100 31.310 41.360 31.570 ;
        RECT 42.010 31.310 42.270 31.570 ;
        RECT 45.210 31.310 45.470 31.570 ;
        RECT 46.850 31.310 47.110 31.570 ;
        RECT 47.760 31.310 48.020 31.570 ;
        RECT 50.960 31.310 51.220 31.570 ;
        RECT 52.600 31.310 52.860 31.570 ;
        RECT 53.510 31.310 53.770 31.570 ;
        RECT 56.710 31.310 56.970 31.570 ;
        RECT 58.350 31.310 58.610 31.570 ;
        RECT 59.260 31.310 59.520 31.570 ;
        RECT 62.460 31.310 62.720 31.570 ;
        RECT 64.100 31.310 64.360 31.570 ;
        RECT 65.010 31.310 65.270 31.570 ;
        RECT 68.210 31.310 68.470 31.570 ;
        RECT 69.850 31.310 70.110 31.570 ;
        RECT 70.760 31.310 71.020 31.570 ;
        RECT 73.960 31.310 74.220 31.570 ;
        RECT 75.600 31.310 75.860 31.570 ;
        RECT 76.510 31.310 76.770 31.570 ;
        RECT 79.710 31.310 79.970 31.570 ;
        RECT 81.350 31.310 81.610 31.570 ;
        RECT 82.260 31.310 82.520 31.570 ;
        RECT 85.460 31.310 85.720 31.570 ;
        RECT 87.100 31.310 87.360 31.570 ;
        RECT 88.010 31.310 88.270 31.570 ;
        RECT 91.210 31.310 91.470 31.570 ;
        RECT 92.850 31.310 93.110 31.570 ;
        RECT 93.760 31.310 94.020 31.570 ;
        RECT 2.990 30.580 3.250 30.840 ;
        RECT 3.900 30.580 4.160 30.840 ;
        RECT 5.540 30.490 5.800 30.750 ;
        RECT 8.740 30.580 9.000 30.840 ;
        RECT 9.650 30.580 9.910 30.840 ;
        RECT 11.290 30.490 11.550 30.750 ;
        RECT 14.490 30.580 14.750 30.840 ;
        RECT 15.400 30.580 15.660 30.840 ;
        RECT 17.040 30.490 17.300 30.750 ;
        RECT 20.240 30.580 20.500 30.840 ;
        RECT 21.150 30.580 21.410 30.840 ;
        RECT 22.790 30.490 23.050 30.750 ;
        RECT 25.990 30.580 26.250 30.840 ;
        RECT 26.900 30.580 27.160 30.840 ;
        RECT 28.540 30.490 28.800 30.750 ;
        RECT 31.740 30.580 32.000 30.840 ;
        RECT 32.650 30.580 32.910 30.840 ;
        RECT 34.290 30.490 34.550 30.750 ;
        RECT 37.490 30.580 37.750 30.840 ;
        RECT 38.400 30.580 38.660 30.840 ;
        RECT 40.040 30.490 40.300 30.750 ;
        RECT 43.240 30.580 43.500 30.840 ;
        RECT 44.150 30.580 44.410 30.840 ;
        RECT 45.790 30.490 46.050 30.750 ;
        RECT 48.990 30.580 49.250 30.840 ;
        RECT 49.900 30.580 50.160 30.840 ;
        RECT 51.540 30.490 51.800 30.750 ;
        RECT 54.740 30.580 55.000 30.840 ;
        RECT 55.650 30.580 55.910 30.840 ;
        RECT 57.290 30.490 57.550 30.750 ;
        RECT 60.490 30.580 60.750 30.840 ;
        RECT 61.400 30.580 61.660 30.840 ;
        RECT 63.040 30.490 63.300 30.750 ;
        RECT 66.240 30.580 66.500 30.840 ;
        RECT 67.150 30.580 67.410 30.840 ;
        RECT 68.790 30.490 69.050 30.750 ;
        RECT 71.990 30.580 72.250 30.840 ;
        RECT 72.900 30.580 73.160 30.840 ;
        RECT 74.540 30.490 74.800 30.750 ;
        RECT 77.740 30.580 78.000 30.840 ;
        RECT 78.650 30.580 78.910 30.840 ;
        RECT 80.290 30.490 80.550 30.750 ;
        RECT 83.490 30.580 83.750 30.840 ;
        RECT 84.400 30.580 84.660 30.840 ;
        RECT 86.040 30.490 86.300 30.750 ;
        RECT 89.240 30.580 89.500 30.840 ;
        RECT 90.150 30.580 90.410 30.840 ;
        RECT 91.790 30.490 92.050 30.750 ;
        RECT 1.290 28.540 1.550 28.800 ;
        RECT 4.960 28.900 5.220 29.160 ;
        RECT 6.600 28.900 6.860 29.160 ;
        RECT 7.510 28.900 7.770 29.160 ;
        RECT 10.710 28.900 10.970 29.160 ;
        RECT 12.350 28.900 12.610 29.160 ;
        RECT 13.260 28.900 13.520 29.160 ;
        RECT 16.460 28.900 16.720 29.160 ;
        RECT 18.100 28.900 18.360 29.160 ;
        RECT 19.010 28.900 19.270 29.160 ;
        RECT 22.210 28.900 22.470 29.160 ;
        RECT 23.850 28.900 24.110 29.160 ;
        RECT 24.760 28.900 25.020 29.160 ;
        RECT 27.960 28.900 28.220 29.160 ;
        RECT 29.600 28.900 29.860 29.160 ;
        RECT 30.510 28.900 30.770 29.160 ;
        RECT 33.710 28.900 33.970 29.160 ;
        RECT 35.350 28.900 35.610 29.160 ;
        RECT 36.260 28.900 36.520 29.160 ;
        RECT 39.460 28.900 39.720 29.160 ;
        RECT 41.100 28.900 41.360 29.160 ;
        RECT 42.010 28.900 42.270 29.160 ;
        RECT 45.210 28.900 45.470 29.160 ;
        RECT 46.850 28.900 47.110 29.160 ;
        RECT 47.760 28.900 48.020 29.160 ;
        RECT 50.960 28.900 51.220 29.160 ;
        RECT 52.600 28.900 52.860 29.160 ;
        RECT 53.510 28.900 53.770 29.160 ;
        RECT 56.710 28.900 56.970 29.160 ;
        RECT 58.350 28.900 58.610 29.160 ;
        RECT 59.260 28.900 59.520 29.160 ;
        RECT 62.460 28.900 62.720 29.160 ;
        RECT 64.100 28.900 64.360 29.160 ;
        RECT 65.010 28.900 65.270 29.160 ;
        RECT 68.210 28.900 68.470 29.160 ;
        RECT 69.850 28.900 70.110 29.160 ;
        RECT 70.760 28.900 71.020 29.160 ;
        RECT 73.960 28.900 74.220 29.160 ;
        RECT 75.600 28.900 75.860 29.160 ;
        RECT 76.510 28.900 76.770 29.160 ;
        RECT 79.710 28.900 79.970 29.160 ;
        RECT 81.350 28.900 81.610 29.160 ;
        RECT 82.260 28.900 82.520 29.160 ;
        RECT 85.460 28.900 85.720 29.160 ;
        RECT 87.100 28.900 87.360 29.160 ;
        RECT 88.010 28.900 88.270 29.160 ;
        RECT 91.210 28.900 91.470 29.160 ;
        RECT 92.850 28.900 93.110 29.160 ;
        RECT 93.760 28.900 94.020 29.160 ;
        RECT 2.990 27.770 3.250 28.030 ;
        RECT 3.900 27.770 4.160 28.030 ;
        RECT 5.540 27.680 5.800 27.940 ;
        RECT 8.740 27.770 9.000 28.030 ;
        RECT 9.650 27.770 9.910 28.030 ;
        RECT 11.290 27.680 11.550 27.940 ;
        RECT 14.490 27.770 14.750 28.030 ;
        RECT 15.400 27.770 15.660 28.030 ;
        RECT 17.040 27.680 17.300 27.940 ;
        RECT 20.240 27.770 20.500 28.030 ;
        RECT 21.150 27.770 21.410 28.030 ;
        RECT 22.790 27.680 23.050 27.940 ;
        RECT 25.990 27.770 26.250 28.030 ;
        RECT 26.900 27.770 27.160 28.030 ;
        RECT 28.540 27.680 28.800 27.940 ;
        RECT 31.740 27.770 32.000 28.030 ;
        RECT 32.650 27.770 32.910 28.030 ;
        RECT 34.290 27.680 34.550 27.940 ;
        RECT 37.490 27.770 37.750 28.030 ;
        RECT 38.400 27.770 38.660 28.030 ;
        RECT 40.040 27.680 40.300 27.940 ;
        RECT 43.240 27.770 43.500 28.030 ;
        RECT 44.150 27.770 44.410 28.030 ;
        RECT 45.790 27.680 46.050 27.940 ;
        RECT 48.990 27.770 49.250 28.030 ;
        RECT 49.900 27.770 50.160 28.030 ;
        RECT 51.540 27.680 51.800 27.940 ;
        RECT 54.740 27.770 55.000 28.030 ;
        RECT 55.650 27.770 55.910 28.030 ;
        RECT 57.290 27.680 57.550 27.940 ;
        RECT 60.490 27.770 60.750 28.030 ;
        RECT 61.400 27.770 61.660 28.030 ;
        RECT 63.040 27.680 63.300 27.940 ;
        RECT 66.240 27.770 66.500 28.030 ;
        RECT 67.150 27.770 67.410 28.030 ;
        RECT 68.790 27.680 69.050 27.940 ;
        RECT 71.990 27.770 72.250 28.030 ;
        RECT 72.900 27.770 73.160 28.030 ;
        RECT 74.540 27.680 74.800 27.940 ;
        RECT 77.740 27.770 78.000 28.030 ;
        RECT 78.650 27.770 78.910 28.030 ;
        RECT 80.290 27.680 80.550 27.940 ;
        RECT 83.490 27.770 83.750 28.030 ;
        RECT 84.400 27.770 84.660 28.030 ;
        RECT 86.040 27.680 86.300 27.940 ;
        RECT 89.240 27.770 89.500 28.030 ;
        RECT 90.150 27.770 90.410 28.030 ;
        RECT 91.790 27.680 92.050 27.940 ;
        RECT 1.280 25.730 1.540 25.990 ;
        RECT 4.960 26.090 5.220 26.350 ;
        RECT 6.600 26.090 6.860 26.350 ;
        RECT 7.510 26.090 7.770 26.350 ;
        RECT 10.710 26.090 10.970 26.350 ;
        RECT 12.350 26.090 12.610 26.350 ;
        RECT 13.260 26.090 13.520 26.350 ;
        RECT 16.460 26.090 16.720 26.350 ;
        RECT 18.100 26.090 18.360 26.350 ;
        RECT 19.010 26.090 19.270 26.350 ;
        RECT 22.210 26.090 22.470 26.350 ;
        RECT 23.850 26.090 24.110 26.350 ;
        RECT 24.760 26.090 25.020 26.350 ;
        RECT 27.960 26.090 28.220 26.350 ;
        RECT 29.600 26.090 29.860 26.350 ;
        RECT 30.510 26.090 30.770 26.350 ;
        RECT 33.710 26.090 33.970 26.350 ;
        RECT 35.350 26.090 35.610 26.350 ;
        RECT 36.260 26.090 36.520 26.350 ;
        RECT 39.460 26.090 39.720 26.350 ;
        RECT 41.100 26.090 41.360 26.350 ;
        RECT 42.010 26.090 42.270 26.350 ;
        RECT 45.210 26.090 45.470 26.350 ;
        RECT 46.850 26.090 47.110 26.350 ;
        RECT 47.760 26.090 48.020 26.350 ;
        RECT 50.960 26.090 51.220 26.350 ;
        RECT 52.600 26.090 52.860 26.350 ;
        RECT 53.510 26.090 53.770 26.350 ;
        RECT 56.710 26.090 56.970 26.350 ;
        RECT 58.350 26.090 58.610 26.350 ;
        RECT 59.260 26.090 59.520 26.350 ;
        RECT 62.460 26.090 62.720 26.350 ;
        RECT 64.100 26.090 64.360 26.350 ;
        RECT 65.010 26.090 65.270 26.350 ;
        RECT 68.210 26.090 68.470 26.350 ;
        RECT 69.850 26.090 70.110 26.350 ;
        RECT 70.760 26.090 71.020 26.350 ;
        RECT 73.960 26.090 74.220 26.350 ;
        RECT 75.600 26.090 75.860 26.350 ;
        RECT 76.510 26.090 76.770 26.350 ;
        RECT 79.710 26.090 79.970 26.350 ;
        RECT 81.350 26.090 81.610 26.350 ;
        RECT 82.260 26.090 82.520 26.350 ;
        RECT 85.460 26.090 85.720 26.350 ;
        RECT 87.100 26.090 87.360 26.350 ;
        RECT 88.010 26.090 88.270 26.350 ;
        RECT 91.210 26.090 91.470 26.350 ;
        RECT 92.850 26.090 93.110 26.350 ;
        RECT 93.760 26.090 94.020 26.350 ;
        RECT 2.990 25.360 3.250 25.620 ;
        RECT 3.900 25.360 4.160 25.620 ;
        RECT 5.540 25.270 5.800 25.530 ;
        RECT 8.740 25.360 9.000 25.620 ;
        RECT 9.650 25.360 9.910 25.620 ;
        RECT 11.290 25.270 11.550 25.530 ;
        RECT 14.490 25.360 14.750 25.620 ;
        RECT 15.400 25.360 15.660 25.620 ;
        RECT 17.040 25.270 17.300 25.530 ;
        RECT 20.240 25.360 20.500 25.620 ;
        RECT 21.150 25.360 21.410 25.620 ;
        RECT 22.790 25.270 23.050 25.530 ;
        RECT 25.990 25.360 26.250 25.620 ;
        RECT 26.900 25.360 27.160 25.620 ;
        RECT 28.540 25.270 28.800 25.530 ;
        RECT 31.740 25.360 32.000 25.620 ;
        RECT 32.650 25.360 32.910 25.620 ;
        RECT 34.290 25.270 34.550 25.530 ;
        RECT 37.490 25.360 37.750 25.620 ;
        RECT 38.400 25.360 38.660 25.620 ;
        RECT 40.040 25.270 40.300 25.530 ;
        RECT 43.240 25.360 43.500 25.620 ;
        RECT 44.150 25.360 44.410 25.620 ;
        RECT 45.790 25.270 46.050 25.530 ;
        RECT 48.990 25.360 49.250 25.620 ;
        RECT 49.900 25.360 50.160 25.620 ;
        RECT 51.540 25.270 51.800 25.530 ;
        RECT 54.740 25.360 55.000 25.620 ;
        RECT 55.650 25.360 55.910 25.620 ;
        RECT 57.290 25.270 57.550 25.530 ;
        RECT 60.490 25.360 60.750 25.620 ;
        RECT 61.400 25.360 61.660 25.620 ;
        RECT 63.040 25.270 63.300 25.530 ;
        RECT 66.240 25.360 66.500 25.620 ;
        RECT 67.150 25.360 67.410 25.620 ;
        RECT 68.790 25.270 69.050 25.530 ;
        RECT 71.990 25.360 72.250 25.620 ;
        RECT 72.900 25.360 73.160 25.620 ;
        RECT 74.540 25.270 74.800 25.530 ;
        RECT 77.740 25.360 78.000 25.620 ;
        RECT 78.650 25.360 78.910 25.620 ;
        RECT 80.290 25.270 80.550 25.530 ;
        RECT 83.490 25.360 83.750 25.620 ;
        RECT 84.400 25.360 84.660 25.620 ;
        RECT 86.040 25.270 86.300 25.530 ;
        RECT 89.240 25.360 89.500 25.620 ;
        RECT 90.150 25.360 90.410 25.620 ;
        RECT 91.790 25.270 92.050 25.530 ;
        RECT 1.290 23.320 1.550 23.580 ;
        RECT 4.960 23.680 5.220 23.940 ;
        RECT 6.600 23.680 6.860 23.940 ;
        RECT 7.510 23.680 7.770 23.940 ;
        RECT 10.710 23.680 10.970 23.940 ;
        RECT 12.350 23.680 12.610 23.940 ;
        RECT 13.260 23.680 13.520 23.940 ;
        RECT 16.460 23.680 16.720 23.940 ;
        RECT 18.100 23.680 18.360 23.940 ;
        RECT 19.010 23.680 19.270 23.940 ;
        RECT 22.210 23.680 22.470 23.940 ;
        RECT 23.850 23.680 24.110 23.940 ;
        RECT 24.760 23.680 25.020 23.940 ;
        RECT 27.960 23.680 28.220 23.940 ;
        RECT 29.600 23.680 29.860 23.940 ;
        RECT 30.510 23.680 30.770 23.940 ;
        RECT 33.710 23.680 33.970 23.940 ;
        RECT 35.350 23.680 35.610 23.940 ;
        RECT 36.260 23.680 36.520 23.940 ;
        RECT 39.460 23.680 39.720 23.940 ;
        RECT 41.100 23.680 41.360 23.940 ;
        RECT 42.010 23.680 42.270 23.940 ;
        RECT 45.210 23.680 45.470 23.940 ;
        RECT 46.850 23.680 47.110 23.940 ;
        RECT 47.760 23.680 48.020 23.940 ;
        RECT 50.960 23.680 51.220 23.940 ;
        RECT 52.600 23.680 52.860 23.940 ;
        RECT 53.510 23.680 53.770 23.940 ;
        RECT 56.710 23.680 56.970 23.940 ;
        RECT 58.350 23.680 58.610 23.940 ;
        RECT 59.260 23.680 59.520 23.940 ;
        RECT 62.460 23.680 62.720 23.940 ;
        RECT 64.100 23.680 64.360 23.940 ;
        RECT 65.010 23.680 65.270 23.940 ;
        RECT 68.210 23.680 68.470 23.940 ;
        RECT 69.850 23.680 70.110 23.940 ;
        RECT 70.760 23.680 71.020 23.940 ;
        RECT 73.960 23.680 74.220 23.940 ;
        RECT 75.600 23.680 75.860 23.940 ;
        RECT 76.510 23.680 76.770 23.940 ;
        RECT 79.710 23.680 79.970 23.940 ;
        RECT 81.350 23.680 81.610 23.940 ;
        RECT 82.260 23.680 82.520 23.940 ;
        RECT 85.460 23.680 85.720 23.940 ;
        RECT 87.100 23.680 87.360 23.940 ;
        RECT 88.010 23.680 88.270 23.940 ;
        RECT 91.210 23.680 91.470 23.940 ;
        RECT 92.850 23.680 93.110 23.940 ;
        RECT 93.760 23.680 94.020 23.940 ;
        RECT 2.990 22.950 3.250 23.210 ;
        RECT 3.900 22.950 4.160 23.210 ;
        RECT 5.540 22.860 5.800 23.120 ;
        RECT 8.740 22.950 9.000 23.210 ;
        RECT 9.650 22.950 9.910 23.210 ;
        RECT 11.290 22.860 11.550 23.120 ;
        RECT 14.490 22.950 14.750 23.210 ;
        RECT 15.400 22.950 15.660 23.210 ;
        RECT 17.040 22.860 17.300 23.120 ;
        RECT 20.240 22.950 20.500 23.210 ;
        RECT 21.150 22.950 21.410 23.210 ;
        RECT 22.790 22.860 23.050 23.120 ;
        RECT 25.990 22.950 26.250 23.210 ;
        RECT 26.900 22.950 27.160 23.210 ;
        RECT 28.540 22.860 28.800 23.120 ;
        RECT 31.740 22.950 32.000 23.210 ;
        RECT 32.650 22.950 32.910 23.210 ;
        RECT 34.290 22.860 34.550 23.120 ;
        RECT 37.490 22.950 37.750 23.210 ;
        RECT 38.400 22.950 38.660 23.210 ;
        RECT 40.040 22.860 40.300 23.120 ;
        RECT 43.240 22.950 43.500 23.210 ;
        RECT 44.150 22.950 44.410 23.210 ;
        RECT 45.790 22.860 46.050 23.120 ;
        RECT 48.990 22.950 49.250 23.210 ;
        RECT 49.900 22.950 50.160 23.210 ;
        RECT 51.540 22.860 51.800 23.120 ;
        RECT 54.740 22.950 55.000 23.210 ;
        RECT 55.650 22.950 55.910 23.210 ;
        RECT 57.290 22.860 57.550 23.120 ;
        RECT 60.490 22.950 60.750 23.210 ;
        RECT 61.400 22.950 61.660 23.210 ;
        RECT 63.040 22.860 63.300 23.120 ;
        RECT 66.240 22.950 66.500 23.210 ;
        RECT 67.150 22.950 67.410 23.210 ;
        RECT 68.790 22.860 69.050 23.120 ;
        RECT 71.990 22.950 72.250 23.210 ;
        RECT 72.900 22.950 73.160 23.210 ;
        RECT 74.540 22.860 74.800 23.120 ;
        RECT 77.740 22.950 78.000 23.210 ;
        RECT 78.650 22.950 78.910 23.210 ;
        RECT 80.290 22.860 80.550 23.120 ;
        RECT 83.490 22.950 83.750 23.210 ;
        RECT 84.400 22.950 84.660 23.210 ;
        RECT 86.040 22.860 86.300 23.120 ;
        RECT 89.240 22.950 89.500 23.210 ;
        RECT 90.150 22.950 90.410 23.210 ;
        RECT 91.790 22.860 92.050 23.120 ;
        RECT 1.290 20.910 1.550 21.170 ;
        RECT 4.960 21.270 5.220 21.530 ;
        RECT 6.600 21.270 6.860 21.530 ;
        RECT 7.510 21.270 7.770 21.530 ;
        RECT 10.710 21.270 10.970 21.530 ;
        RECT 12.350 21.270 12.610 21.530 ;
        RECT 13.260 21.270 13.520 21.530 ;
        RECT 16.460 21.270 16.720 21.530 ;
        RECT 18.100 21.270 18.360 21.530 ;
        RECT 19.010 21.270 19.270 21.530 ;
        RECT 22.210 21.270 22.470 21.530 ;
        RECT 23.850 21.270 24.110 21.530 ;
        RECT 24.760 21.270 25.020 21.530 ;
        RECT 27.960 21.270 28.220 21.530 ;
        RECT 29.600 21.270 29.860 21.530 ;
        RECT 30.510 21.270 30.770 21.530 ;
        RECT 33.710 21.270 33.970 21.530 ;
        RECT 35.350 21.270 35.610 21.530 ;
        RECT 36.260 21.270 36.520 21.530 ;
        RECT 39.460 21.270 39.720 21.530 ;
        RECT 41.100 21.270 41.360 21.530 ;
        RECT 42.010 21.270 42.270 21.530 ;
        RECT 45.210 21.270 45.470 21.530 ;
        RECT 46.850 21.270 47.110 21.530 ;
        RECT 47.760 21.270 48.020 21.530 ;
        RECT 50.960 21.270 51.220 21.530 ;
        RECT 52.600 21.270 52.860 21.530 ;
        RECT 53.510 21.270 53.770 21.530 ;
        RECT 56.710 21.270 56.970 21.530 ;
        RECT 58.350 21.270 58.610 21.530 ;
        RECT 59.260 21.270 59.520 21.530 ;
        RECT 62.460 21.270 62.720 21.530 ;
        RECT 64.100 21.270 64.360 21.530 ;
        RECT 65.010 21.270 65.270 21.530 ;
        RECT 68.210 21.270 68.470 21.530 ;
        RECT 69.850 21.270 70.110 21.530 ;
        RECT 70.760 21.270 71.020 21.530 ;
        RECT 73.960 21.270 74.220 21.530 ;
        RECT 75.600 21.270 75.860 21.530 ;
        RECT 76.510 21.270 76.770 21.530 ;
        RECT 79.710 21.270 79.970 21.530 ;
        RECT 81.350 21.270 81.610 21.530 ;
        RECT 82.260 21.270 82.520 21.530 ;
        RECT 85.460 21.270 85.720 21.530 ;
        RECT 87.100 21.270 87.360 21.530 ;
        RECT 88.010 21.270 88.270 21.530 ;
        RECT 91.210 21.270 91.470 21.530 ;
        RECT 92.850 21.270 93.110 21.530 ;
        RECT 93.760 21.270 94.020 21.530 ;
        RECT 2.990 20.540 3.250 20.800 ;
        RECT 3.900 20.540 4.160 20.800 ;
        RECT 5.540 20.450 5.800 20.710 ;
        RECT 8.740 20.540 9.000 20.800 ;
        RECT 9.650 20.540 9.910 20.800 ;
        RECT 11.290 20.450 11.550 20.710 ;
        RECT 14.490 20.540 14.750 20.800 ;
        RECT 15.400 20.540 15.660 20.800 ;
        RECT 17.040 20.450 17.300 20.710 ;
        RECT 20.240 20.540 20.500 20.800 ;
        RECT 21.150 20.540 21.410 20.800 ;
        RECT 22.790 20.450 23.050 20.710 ;
        RECT 25.990 20.540 26.250 20.800 ;
        RECT 26.900 20.540 27.160 20.800 ;
        RECT 28.540 20.450 28.800 20.710 ;
        RECT 31.740 20.540 32.000 20.800 ;
        RECT 32.650 20.540 32.910 20.800 ;
        RECT 34.290 20.450 34.550 20.710 ;
        RECT 37.490 20.540 37.750 20.800 ;
        RECT 38.400 20.540 38.660 20.800 ;
        RECT 40.040 20.450 40.300 20.710 ;
        RECT 43.240 20.540 43.500 20.800 ;
        RECT 44.150 20.540 44.410 20.800 ;
        RECT 45.790 20.450 46.050 20.710 ;
        RECT 48.990 20.540 49.250 20.800 ;
        RECT 49.900 20.540 50.160 20.800 ;
        RECT 51.540 20.450 51.800 20.710 ;
        RECT 54.740 20.540 55.000 20.800 ;
        RECT 55.650 20.540 55.910 20.800 ;
        RECT 57.290 20.450 57.550 20.710 ;
        RECT 60.490 20.540 60.750 20.800 ;
        RECT 61.400 20.540 61.660 20.800 ;
        RECT 63.040 20.450 63.300 20.710 ;
        RECT 66.240 20.540 66.500 20.800 ;
        RECT 67.150 20.540 67.410 20.800 ;
        RECT 68.790 20.450 69.050 20.710 ;
        RECT 71.990 20.540 72.250 20.800 ;
        RECT 72.900 20.540 73.160 20.800 ;
        RECT 74.540 20.450 74.800 20.710 ;
        RECT 77.740 20.540 78.000 20.800 ;
        RECT 78.650 20.540 78.910 20.800 ;
        RECT 80.290 20.450 80.550 20.710 ;
        RECT 83.490 20.540 83.750 20.800 ;
        RECT 84.400 20.540 84.660 20.800 ;
        RECT 86.040 20.450 86.300 20.710 ;
        RECT 89.240 20.540 89.500 20.800 ;
        RECT 90.150 20.540 90.410 20.800 ;
        RECT 91.790 20.450 92.050 20.710 ;
        RECT 1.290 18.500 1.550 18.760 ;
        RECT 4.960 18.860 5.220 19.120 ;
        RECT 6.600 18.860 6.860 19.120 ;
        RECT 7.510 18.860 7.770 19.120 ;
        RECT 10.710 18.860 10.970 19.120 ;
        RECT 12.350 18.860 12.610 19.120 ;
        RECT 13.260 18.860 13.520 19.120 ;
        RECT 16.460 18.860 16.720 19.120 ;
        RECT 18.100 18.860 18.360 19.120 ;
        RECT 19.010 18.860 19.270 19.120 ;
        RECT 22.210 18.860 22.470 19.120 ;
        RECT 23.850 18.860 24.110 19.120 ;
        RECT 24.760 18.860 25.020 19.120 ;
        RECT 27.960 18.860 28.220 19.120 ;
        RECT 29.600 18.860 29.860 19.120 ;
        RECT 30.510 18.860 30.770 19.120 ;
        RECT 33.710 18.860 33.970 19.120 ;
        RECT 35.350 18.860 35.610 19.120 ;
        RECT 36.260 18.860 36.520 19.120 ;
        RECT 39.460 18.860 39.720 19.120 ;
        RECT 41.100 18.860 41.360 19.120 ;
        RECT 42.010 18.860 42.270 19.120 ;
        RECT 45.210 18.860 45.470 19.120 ;
        RECT 46.850 18.860 47.110 19.120 ;
        RECT 47.760 18.860 48.020 19.120 ;
        RECT 50.960 18.860 51.220 19.120 ;
        RECT 52.600 18.860 52.860 19.120 ;
        RECT 53.510 18.860 53.770 19.120 ;
        RECT 56.710 18.860 56.970 19.120 ;
        RECT 58.350 18.860 58.610 19.120 ;
        RECT 59.260 18.860 59.520 19.120 ;
        RECT 62.460 18.860 62.720 19.120 ;
        RECT 64.100 18.860 64.360 19.120 ;
        RECT 65.010 18.860 65.270 19.120 ;
        RECT 68.210 18.860 68.470 19.120 ;
        RECT 69.850 18.860 70.110 19.120 ;
        RECT 70.760 18.860 71.020 19.120 ;
        RECT 73.960 18.860 74.220 19.120 ;
        RECT 75.600 18.860 75.860 19.120 ;
        RECT 76.510 18.860 76.770 19.120 ;
        RECT 79.710 18.860 79.970 19.120 ;
        RECT 81.350 18.860 81.610 19.120 ;
        RECT 82.260 18.860 82.520 19.120 ;
        RECT 85.460 18.860 85.720 19.120 ;
        RECT 87.100 18.860 87.360 19.120 ;
        RECT 88.010 18.860 88.270 19.120 ;
        RECT 91.210 18.860 91.470 19.120 ;
        RECT 92.850 18.860 93.110 19.120 ;
        RECT 93.760 18.860 94.020 19.120 ;
        RECT 2.990 18.130 3.250 18.390 ;
        RECT 3.900 18.130 4.160 18.390 ;
        RECT 5.540 18.040 5.800 18.300 ;
        RECT 8.740 18.130 9.000 18.390 ;
        RECT 9.650 18.130 9.910 18.390 ;
        RECT 11.290 18.040 11.550 18.300 ;
        RECT 14.490 18.130 14.750 18.390 ;
        RECT 15.400 18.130 15.660 18.390 ;
        RECT 17.040 18.040 17.300 18.300 ;
        RECT 20.240 18.130 20.500 18.390 ;
        RECT 21.150 18.130 21.410 18.390 ;
        RECT 22.790 18.040 23.050 18.300 ;
        RECT 25.990 18.130 26.250 18.390 ;
        RECT 26.900 18.130 27.160 18.390 ;
        RECT 28.540 18.040 28.800 18.300 ;
        RECT 31.740 18.130 32.000 18.390 ;
        RECT 32.650 18.130 32.910 18.390 ;
        RECT 34.290 18.040 34.550 18.300 ;
        RECT 37.490 18.130 37.750 18.390 ;
        RECT 38.400 18.130 38.660 18.390 ;
        RECT 40.040 18.040 40.300 18.300 ;
        RECT 43.240 18.130 43.500 18.390 ;
        RECT 44.150 18.130 44.410 18.390 ;
        RECT 45.790 18.040 46.050 18.300 ;
        RECT 48.990 18.130 49.250 18.390 ;
        RECT 49.900 18.130 50.160 18.390 ;
        RECT 51.540 18.040 51.800 18.300 ;
        RECT 54.740 18.130 55.000 18.390 ;
        RECT 55.650 18.130 55.910 18.390 ;
        RECT 57.290 18.040 57.550 18.300 ;
        RECT 60.490 18.130 60.750 18.390 ;
        RECT 61.400 18.130 61.660 18.390 ;
        RECT 63.040 18.040 63.300 18.300 ;
        RECT 66.240 18.130 66.500 18.390 ;
        RECT 67.150 18.130 67.410 18.390 ;
        RECT 68.790 18.040 69.050 18.300 ;
        RECT 71.990 18.130 72.250 18.390 ;
        RECT 72.900 18.130 73.160 18.390 ;
        RECT 74.540 18.040 74.800 18.300 ;
        RECT 77.740 18.130 78.000 18.390 ;
        RECT 78.650 18.130 78.910 18.390 ;
        RECT 80.290 18.040 80.550 18.300 ;
        RECT 83.490 18.130 83.750 18.390 ;
        RECT 84.400 18.130 84.660 18.390 ;
        RECT 86.040 18.040 86.300 18.300 ;
        RECT 89.240 18.130 89.500 18.390 ;
        RECT 90.150 18.130 90.410 18.390 ;
        RECT 91.790 18.040 92.050 18.300 ;
        RECT 1.290 16.090 1.550 16.350 ;
        RECT 4.960 16.450 5.220 16.710 ;
        RECT 6.600 16.450 6.860 16.710 ;
        RECT 7.510 16.450 7.770 16.710 ;
        RECT 10.710 16.450 10.970 16.710 ;
        RECT 12.350 16.450 12.610 16.710 ;
        RECT 13.260 16.450 13.520 16.710 ;
        RECT 16.460 16.450 16.720 16.710 ;
        RECT 18.100 16.450 18.360 16.710 ;
        RECT 19.010 16.450 19.270 16.710 ;
        RECT 22.210 16.450 22.470 16.710 ;
        RECT 23.850 16.450 24.110 16.710 ;
        RECT 24.760 16.450 25.020 16.710 ;
        RECT 27.960 16.450 28.220 16.710 ;
        RECT 29.600 16.450 29.860 16.710 ;
        RECT 30.510 16.450 30.770 16.710 ;
        RECT 33.710 16.450 33.970 16.710 ;
        RECT 35.350 16.450 35.610 16.710 ;
        RECT 36.260 16.450 36.520 16.710 ;
        RECT 39.460 16.450 39.720 16.710 ;
        RECT 41.100 16.450 41.360 16.710 ;
        RECT 42.010 16.450 42.270 16.710 ;
        RECT 45.210 16.450 45.470 16.710 ;
        RECT 46.850 16.450 47.110 16.710 ;
        RECT 47.760 16.450 48.020 16.710 ;
        RECT 50.960 16.450 51.220 16.710 ;
        RECT 52.600 16.450 52.860 16.710 ;
        RECT 53.510 16.450 53.770 16.710 ;
        RECT 56.710 16.450 56.970 16.710 ;
        RECT 58.350 16.450 58.610 16.710 ;
        RECT 59.260 16.450 59.520 16.710 ;
        RECT 62.460 16.450 62.720 16.710 ;
        RECT 64.100 16.450 64.360 16.710 ;
        RECT 65.010 16.450 65.270 16.710 ;
        RECT 68.210 16.450 68.470 16.710 ;
        RECT 69.850 16.450 70.110 16.710 ;
        RECT 70.760 16.450 71.020 16.710 ;
        RECT 73.960 16.450 74.220 16.710 ;
        RECT 75.600 16.450 75.860 16.710 ;
        RECT 76.510 16.450 76.770 16.710 ;
        RECT 79.710 16.450 79.970 16.710 ;
        RECT 81.350 16.450 81.610 16.710 ;
        RECT 82.260 16.450 82.520 16.710 ;
        RECT 85.460 16.450 85.720 16.710 ;
        RECT 87.100 16.450 87.360 16.710 ;
        RECT 88.010 16.450 88.270 16.710 ;
        RECT 91.210 16.450 91.470 16.710 ;
        RECT 92.850 16.450 93.110 16.710 ;
        RECT 93.760 16.450 94.020 16.710 ;
        RECT 2.990 15.720 3.250 15.980 ;
        RECT 3.900 15.720 4.160 15.980 ;
        RECT 5.540 15.630 5.800 15.890 ;
        RECT 8.740 15.720 9.000 15.980 ;
        RECT 9.650 15.720 9.910 15.980 ;
        RECT 11.290 15.630 11.550 15.890 ;
        RECT 14.490 15.720 14.750 15.980 ;
        RECT 15.400 15.720 15.660 15.980 ;
        RECT 17.040 15.630 17.300 15.890 ;
        RECT 20.240 15.720 20.500 15.980 ;
        RECT 21.150 15.720 21.410 15.980 ;
        RECT 22.790 15.630 23.050 15.890 ;
        RECT 25.990 15.720 26.250 15.980 ;
        RECT 26.900 15.720 27.160 15.980 ;
        RECT 28.540 15.630 28.800 15.890 ;
        RECT 31.740 15.720 32.000 15.980 ;
        RECT 32.650 15.720 32.910 15.980 ;
        RECT 34.290 15.630 34.550 15.890 ;
        RECT 37.490 15.720 37.750 15.980 ;
        RECT 38.400 15.720 38.660 15.980 ;
        RECT 40.040 15.630 40.300 15.890 ;
        RECT 43.240 15.720 43.500 15.980 ;
        RECT 44.150 15.720 44.410 15.980 ;
        RECT 45.790 15.630 46.050 15.890 ;
        RECT 48.990 15.720 49.250 15.980 ;
        RECT 49.900 15.720 50.160 15.980 ;
        RECT 51.540 15.630 51.800 15.890 ;
        RECT 54.740 15.720 55.000 15.980 ;
        RECT 55.650 15.720 55.910 15.980 ;
        RECT 57.290 15.630 57.550 15.890 ;
        RECT 60.490 15.720 60.750 15.980 ;
        RECT 61.400 15.720 61.660 15.980 ;
        RECT 63.040 15.630 63.300 15.890 ;
        RECT 66.240 15.720 66.500 15.980 ;
        RECT 67.150 15.720 67.410 15.980 ;
        RECT 68.790 15.630 69.050 15.890 ;
        RECT 71.990 15.720 72.250 15.980 ;
        RECT 72.900 15.720 73.160 15.980 ;
        RECT 74.540 15.630 74.800 15.890 ;
        RECT 77.740 15.720 78.000 15.980 ;
        RECT 78.650 15.720 78.910 15.980 ;
        RECT 80.290 15.630 80.550 15.890 ;
        RECT 83.490 15.720 83.750 15.980 ;
        RECT 84.400 15.720 84.660 15.980 ;
        RECT 86.040 15.630 86.300 15.890 ;
        RECT 89.240 15.720 89.500 15.980 ;
        RECT 90.150 15.720 90.410 15.980 ;
        RECT 91.790 15.630 92.050 15.890 ;
        RECT 1.290 13.680 1.550 13.940 ;
        RECT 4.960 14.040 5.220 14.300 ;
        RECT 6.600 14.040 6.860 14.300 ;
        RECT 7.510 14.040 7.770 14.300 ;
        RECT 10.710 14.040 10.970 14.300 ;
        RECT 12.350 14.040 12.610 14.300 ;
        RECT 13.260 14.040 13.520 14.300 ;
        RECT 16.460 14.040 16.720 14.300 ;
        RECT 18.100 14.040 18.360 14.300 ;
        RECT 19.010 14.040 19.270 14.300 ;
        RECT 22.210 14.040 22.470 14.300 ;
        RECT 23.850 14.040 24.110 14.300 ;
        RECT 24.760 14.040 25.020 14.300 ;
        RECT 27.960 14.040 28.220 14.300 ;
        RECT 29.600 14.040 29.860 14.300 ;
        RECT 30.510 14.040 30.770 14.300 ;
        RECT 33.710 14.040 33.970 14.300 ;
        RECT 35.350 14.040 35.610 14.300 ;
        RECT 36.260 14.040 36.520 14.300 ;
        RECT 39.460 14.040 39.720 14.300 ;
        RECT 41.100 14.040 41.360 14.300 ;
        RECT 42.010 14.040 42.270 14.300 ;
        RECT 45.210 14.040 45.470 14.300 ;
        RECT 46.850 14.040 47.110 14.300 ;
        RECT 47.760 14.040 48.020 14.300 ;
        RECT 50.960 14.040 51.220 14.300 ;
        RECT 52.600 14.040 52.860 14.300 ;
        RECT 53.510 14.040 53.770 14.300 ;
        RECT 56.710 14.040 56.970 14.300 ;
        RECT 58.350 14.040 58.610 14.300 ;
        RECT 59.260 14.040 59.520 14.300 ;
        RECT 62.460 14.040 62.720 14.300 ;
        RECT 64.100 14.040 64.360 14.300 ;
        RECT 65.010 14.040 65.270 14.300 ;
        RECT 68.210 14.040 68.470 14.300 ;
        RECT 69.850 14.040 70.110 14.300 ;
        RECT 70.760 14.040 71.020 14.300 ;
        RECT 73.960 14.040 74.220 14.300 ;
        RECT 75.600 14.040 75.860 14.300 ;
        RECT 76.510 14.040 76.770 14.300 ;
        RECT 79.710 14.040 79.970 14.300 ;
        RECT 81.350 14.040 81.610 14.300 ;
        RECT 82.260 14.040 82.520 14.300 ;
        RECT 85.460 14.040 85.720 14.300 ;
        RECT 87.100 14.040 87.360 14.300 ;
        RECT 88.010 14.040 88.270 14.300 ;
        RECT 91.210 14.040 91.470 14.300 ;
        RECT 92.850 14.040 93.110 14.300 ;
        RECT 93.760 14.040 94.020 14.300 ;
        RECT 2.990 13.310 3.250 13.570 ;
        RECT 3.900 13.310 4.160 13.570 ;
        RECT 5.540 13.220 5.800 13.480 ;
        RECT 8.740 13.310 9.000 13.570 ;
        RECT 9.650 13.310 9.910 13.570 ;
        RECT 11.290 13.220 11.550 13.480 ;
        RECT 14.490 13.310 14.750 13.570 ;
        RECT 15.400 13.310 15.660 13.570 ;
        RECT 17.040 13.220 17.300 13.480 ;
        RECT 20.240 13.310 20.500 13.570 ;
        RECT 21.150 13.310 21.410 13.570 ;
        RECT 22.790 13.220 23.050 13.480 ;
        RECT 25.990 13.310 26.250 13.570 ;
        RECT 26.900 13.310 27.160 13.570 ;
        RECT 28.540 13.220 28.800 13.480 ;
        RECT 31.740 13.310 32.000 13.570 ;
        RECT 32.650 13.310 32.910 13.570 ;
        RECT 34.290 13.220 34.550 13.480 ;
        RECT 37.490 13.310 37.750 13.570 ;
        RECT 38.400 13.310 38.660 13.570 ;
        RECT 40.040 13.220 40.300 13.480 ;
        RECT 43.240 13.310 43.500 13.570 ;
        RECT 44.150 13.310 44.410 13.570 ;
        RECT 45.790 13.220 46.050 13.480 ;
        RECT 48.990 13.310 49.250 13.570 ;
        RECT 49.900 13.310 50.160 13.570 ;
        RECT 51.540 13.220 51.800 13.480 ;
        RECT 54.740 13.310 55.000 13.570 ;
        RECT 55.650 13.310 55.910 13.570 ;
        RECT 57.290 13.220 57.550 13.480 ;
        RECT 60.490 13.310 60.750 13.570 ;
        RECT 61.400 13.310 61.660 13.570 ;
        RECT 63.040 13.220 63.300 13.480 ;
        RECT 66.240 13.310 66.500 13.570 ;
        RECT 67.150 13.310 67.410 13.570 ;
        RECT 68.790 13.220 69.050 13.480 ;
        RECT 71.990 13.310 72.250 13.570 ;
        RECT 72.900 13.310 73.160 13.570 ;
        RECT 74.540 13.220 74.800 13.480 ;
        RECT 77.740 13.310 78.000 13.570 ;
        RECT 78.650 13.310 78.910 13.570 ;
        RECT 80.290 13.220 80.550 13.480 ;
        RECT 83.490 13.310 83.750 13.570 ;
        RECT 84.400 13.310 84.660 13.570 ;
        RECT 86.040 13.220 86.300 13.480 ;
        RECT 89.240 13.310 89.500 13.570 ;
        RECT 90.150 13.310 90.410 13.570 ;
        RECT 91.790 13.220 92.050 13.480 ;
        RECT 1.280 11.270 1.540 11.530 ;
        RECT 4.960 11.630 5.220 11.890 ;
        RECT 6.600 11.630 6.860 11.890 ;
        RECT 7.510 11.630 7.770 11.890 ;
        RECT 10.710 11.630 10.970 11.890 ;
        RECT 12.350 11.630 12.610 11.890 ;
        RECT 13.260 11.630 13.520 11.890 ;
        RECT 16.460 11.630 16.720 11.890 ;
        RECT 18.100 11.630 18.360 11.890 ;
        RECT 19.010 11.630 19.270 11.890 ;
        RECT 22.210 11.630 22.470 11.890 ;
        RECT 23.850 11.630 24.110 11.890 ;
        RECT 24.760 11.630 25.020 11.890 ;
        RECT 27.960 11.630 28.220 11.890 ;
        RECT 29.600 11.630 29.860 11.890 ;
        RECT 30.510 11.630 30.770 11.890 ;
        RECT 33.710 11.630 33.970 11.890 ;
        RECT 35.350 11.630 35.610 11.890 ;
        RECT 36.260 11.630 36.520 11.890 ;
        RECT 39.460 11.630 39.720 11.890 ;
        RECT 41.100 11.630 41.360 11.890 ;
        RECT 42.010 11.630 42.270 11.890 ;
        RECT 45.210 11.630 45.470 11.890 ;
        RECT 46.850 11.630 47.110 11.890 ;
        RECT 47.760 11.630 48.020 11.890 ;
        RECT 50.960 11.630 51.220 11.890 ;
        RECT 52.600 11.630 52.860 11.890 ;
        RECT 53.510 11.630 53.770 11.890 ;
        RECT 56.710 11.630 56.970 11.890 ;
        RECT 58.350 11.630 58.610 11.890 ;
        RECT 59.260 11.630 59.520 11.890 ;
        RECT 62.460 11.630 62.720 11.890 ;
        RECT 64.100 11.630 64.360 11.890 ;
        RECT 65.010 11.630 65.270 11.890 ;
        RECT 68.210 11.630 68.470 11.890 ;
        RECT 69.850 11.630 70.110 11.890 ;
        RECT 70.760 11.630 71.020 11.890 ;
        RECT 73.960 11.630 74.220 11.890 ;
        RECT 75.600 11.630 75.860 11.890 ;
        RECT 76.510 11.630 76.770 11.890 ;
        RECT 79.710 11.630 79.970 11.890 ;
        RECT 81.350 11.630 81.610 11.890 ;
        RECT 82.260 11.630 82.520 11.890 ;
        RECT 85.460 11.630 85.720 11.890 ;
        RECT 87.100 11.630 87.360 11.890 ;
        RECT 88.010 11.630 88.270 11.890 ;
        RECT 91.210 11.630 91.470 11.890 ;
        RECT 92.850 11.630 93.110 11.890 ;
        RECT 93.760 11.630 94.020 11.890 ;
        RECT 2.990 10.900 3.250 11.160 ;
        RECT 3.900 10.900 4.160 11.160 ;
        RECT 5.540 10.810 5.800 11.070 ;
        RECT 8.740 10.900 9.000 11.160 ;
        RECT 9.650 10.900 9.910 11.160 ;
        RECT 11.290 10.810 11.550 11.070 ;
        RECT 14.490 10.900 14.750 11.160 ;
        RECT 15.400 10.900 15.660 11.160 ;
        RECT 17.040 10.810 17.300 11.070 ;
        RECT 20.240 10.900 20.500 11.160 ;
        RECT 21.150 10.900 21.410 11.160 ;
        RECT 22.790 10.810 23.050 11.070 ;
        RECT 25.990 10.900 26.250 11.160 ;
        RECT 26.900 10.900 27.160 11.160 ;
        RECT 28.540 10.810 28.800 11.070 ;
        RECT 31.740 10.900 32.000 11.160 ;
        RECT 32.650 10.900 32.910 11.160 ;
        RECT 34.290 10.810 34.550 11.070 ;
        RECT 37.490 10.900 37.750 11.160 ;
        RECT 38.400 10.900 38.660 11.160 ;
        RECT 40.040 10.810 40.300 11.070 ;
        RECT 43.240 10.900 43.500 11.160 ;
        RECT 44.150 10.900 44.410 11.160 ;
        RECT 45.790 10.810 46.050 11.070 ;
        RECT 48.990 10.900 49.250 11.160 ;
        RECT 49.900 10.900 50.160 11.160 ;
        RECT 51.540 10.810 51.800 11.070 ;
        RECT 54.740 10.900 55.000 11.160 ;
        RECT 55.650 10.900 55.910 11.160 ;
        RECT 57.290 10.810 57.550 11.070 ;
        RECT 60.490 10.900 60.750 11.160 ;
        RECT 61.400 10.900 61.660 11.160 ;
        RECT 63.040 10.810 63.300 11.070 ;
        RECT 66.240 10.900 66.500 11.160 ;
        RECT 67.150 10.900 67.410 11.160 ;
        RECT 68.790 10.810 69.050 11.070 ;
        RECT 71.990 10.900 72.250 11.160 ;
        RECT 72.900 10.900 73.160 11.160 ;
        RECT 74.540 10.810 74.800 11.070 ;
        RECT 77.740 10.900 78.000 11.160 ;
        RECT 78.650 10.900 78.910 11.160 ;
        RECT 80.290 10.810 80.550 11.070 ;
        RECT 83.490 10.900 83.750 11.160 ;
        RECT 84.400 10.900 84.660 11.160 ;
        RECT 86.040 10.810 86.300 11.070 ;
        RECT 89.240 10.900 89.500 11.160 ;
        RECT 90.150 10.900 90.410 11.160 ;
        RECT 91.790 10.810 92.050 11.070 ;
        RECT 1.290 8.860 1.550 9.120 ;
        RECT 4.960 9.220 5.220 9.480 ;
        RECT 6.600 9.220 6.860 9.480 ;
        RECT 7.510 9.220 7.770 9.480 ;
        RECT 10.710 9.220 10.970 9.480 ;
        RECT 12.350 9.220 12.610 9.480 ;
        RECT 13.260 9.220 13.520 9.480 ;
        RECT 16.460 9.220 16.720 9.480 ;
        RECT 18.100 9.220 18.360 9.480 ;
        RECT 19.010 9.220 19.270 9.480 ;
        RECT 22.210 9.220 22.470 9.480 ;
        RECT 23.850 9.220 24.110 9.480 ;
        RECT 24.760 9.220 25.020 9.480 ;
        RECT 27.960 9.220 28.220 9.480 ;
        RECT 29.600 9.220 29.860 9.480 ;
        RECT 30.510 9.220 30.770 9.480 ;
        RECT 33.710 9.220 33.970 9.480 ;
        RECT 35.350 9.220 35.610 9.480 ;
        RECT 36.260 9.220 36.520 9.480 ;
        RECT 39.460 9.220 39.720 9.480 ;
        RECT 41.100 9.220 41.360 9.480 ;
        RECT 42.010 9.220 42.270 9.480 ;
        RECT 45.210 9.220 45.470 9.480 ;
        RECT 46.850 9.220 47.110 9.480 ;
        RECT 47.760 9.220 48.020 9.480 ;
        RECT 50.960 9.220 51.220 9.480 ;
        RECT 52.600 9.220 52.860 9.480 ;
        RECT 53.510 9.220 53.770 9.480 ;
        RECT 56.710 9.220 56.970 9.480 ;
        RECT 58.350 9.220 58.610 9.480 ;
        RECT 59.260 9.220 59.520 9.480 ;
        RECT 62.460 9.220 62.720 9.480 ;
        RECT 64.100 9.220 64.360 9.480 ;
        RECT 65.010 9.220 65.270 9.480 ;
        RECT 68.210 9.220 68.470 9.480 ;
        RECT 69.850 9.220 70.110 9.480 ;
        RECT 70.760 9.220 71.020 9.480 ;
        RECT 73.960 9.220 74.220 9.480 ;
        RECT 75.600 9.220 75.860 9.480 ;
        RECT 76.510 9.220 76.770 9.480 ;
        RECT 79.710 9.220 79.970 9.480 ;
        RECT 81.350 9.220 81.610 9.480 ;
        RECT 82.260 9.220 82.520 9.480 ;
        RECT 85.460 9.220 85.720 9.480 ;
        RECT 87.100 9.220 87.360 9.480 ;
        RECT 88.010 9.220 88.270 9.480 ;
        RECT 91.210 9.220 91.470 9.480 ;
        RECT 92.850 9.220 93.110 9.480 ;
        RECT 93.760 9.220 94.020 9.480 ;
        RECT 2.990 8.080 3.250 8.340 ;
        RECT 3.900 8.080 4.160 8.340 ;
        RECT 5.540 7.990 5.800 8.250 ;
        RECT 8.740 8.080 9.000 8.340 ;
        RECT 9.650 8.080 9.910 8.340 ;
        RECT 11.290 7.990 11.550 8.250 ;
        RECT 14.490 8.080 14.750 8.340 ;
        RECT 15.400 8.080 15.660 8.340 ;
        RECT 17.040 7.990 17.300 8.250 ;
        RECT 20.240 8.080 20.500 8.340 ;
        RECT 21.150 8.080 21.410 8.340 ;
        RECT 22.790 7.990 23.050 8.250 ;
        RECT 25.990 8.080 26.250 8.340 ;
        RECT 26.900 8.080 27.160 8.340 ;
        RECT 28.540 7.990 28.800 8.250 ;
        RECT 31.740 8.080 32.000 8.340 ;
        RECT 32.650 8.080 32.910 8.340 ;
        RECT 34.290 7.990 34.550 8.250 ;
        RECT 37.490 8.080 37.750 8.340 ;
        RECT 38.400 8.080 38.660 8.340 ;
        RECT 40.040 7.990 40.300 8.250 ;
        RECT 43.240 8.080 43.500 8.340 ;
        RECT 44.150 8.080 44.410 8.340 ;
        RECT 45.790 7.990 46.050 8.250 ;
        RECT 48.990 8.080 49.250 8.340 ;
        RECT 49.900 8.080 50.160 8.340 ;
        RECT 51.540 7.990 51.800 8.250 ;
        RECT 54.740 8.080 55.000 8.340 ;
        RECT 55.650 8.080 55.910 8.340 ;
        RECT 57.290 7.990 57.550 8.250 ;
        RECT 60.490 8.080 60.750 8.340 ;
        RECT 61.400 8.080 61.660 8.340 ;
        RECT 63.040 7.990 63.300 8.250 ;
        RECT 66.240 8.080 66.500 8.340 ;
        RECT 67.150 8.080 67.410 8.340 ;
        RECT 68.790 7.990 69.050 8.250 ;
        RECT 71.990 8.080 72.250 8.340 ;
        RECT 72.900 8.080 73.160 8.340 ;
        RECT 74.540 7.990 74.800 8.250 ;
        RECT 77.740 8.080 78.000 8.340 ;
        RECT 78.650 8.080 78.910 8.340 ;
        RECT 80.290 7.990 80.550 8.250 ;
        RECT 83.490 8.080 83.750 8.340 ;
        RECT 84.400 8.080 84.660 8.340 ;
        RECT 86.040 7.990 86.300 8.250 ;
        RECT 89.240 8.080 89.500 8.340 ;
        RECT 90.150 8.080 90.410 8.340 ;
        RECT 91.790 7.990 92.050 8.250 ;
        RECT 1.280 6.040 1.540 6.300 ;
        RECT 4.960 6.400 5.220 6.660 ;
        RECT 6.600 6.400 6.860 6.660 ;
        RECT 7.510 6.400 7.770 6.660 ;
        RECT 10.710 6.400 10.970 6.660 ;
        RECT 12.350 6.400 12.610 6.660 ;
        RECT 13.260 6.400 13.520 6.660 ;
        RECT 16.460 6.400 16.720 6.660 ;
        RECT 18.100 6.400 18.360 6.660 ;
        RECT 19.010 6.400 19.270 6.660 ;
        RECT 22.210 6.400 22.470 6.660 ;
        RECT 23.850 6.400 24.110 6.660 ;
        RECT 24.760 6.400 25.020 6.660 ;
        RECT 27.960 6.400 28.220 6.660 ;
        RECT 29.600 6.400 29.860 6.660 ;
        RECT 30.510 6.400 30.770 6.660 ;
        RECT 33.710 6.400 33.970 6.660 ;
        RECT 35.350 6.400 35.610 6.660 ;
        RECT 36.260 6.400 36.520 6.660 ;
        RECT 39.460 6.400 39.720 6.660 ;
        RECT 41.100 6.400 41.360 6.660 ;
        RECT 42.010 6.400 42.270 6.660 ;
        RECT 45.210 6.400 45.470 6.660 ;
        RECT 46.850 6.400 47.110 6.660 ;
        RECT 47.760 6.400 48.020 6.660 ;
        RECT 50.960 6.400 51.220 6.660 ;
        RECT 52.600 6.400 52.860 6.660 ;
        RECT 53.510 6.400 53.770 6.660 ;
        RECT 56.710 6.400 56.970 6.660 ;
        RECT 58.350 6.400 58.610 6.660 ;
        RECT 59.260 6.400 59.520 6.660 ;
        RECT 62.460 6.400 62.720 6.660 ;
        RECT 64.100 6.400 64.360 6.660 ;
        RECT 65.010 6.400 65.270 6.660 ;
        RECT 68.210 6.400 68.470 6.660 ;
        RECT 69.850 6.400 70.110 6.660 ;
        RECT 70.760 6.400 71.020 6.660 ;
        RECT 73.960 6.400 74.220 6.660 ;
        RECT 75.600 6.400 75.860 6.660 ;
        RECT 76.510 6.400 76.770 6.660 ;
        RECT 79.710 6.400 79.970 6.660 ;
        RECT 81.350 6.400 81.610 6.660 ;
        RECT 82.260 6.400 82.520 6.660 ;
        RECT 85.460 6.400 85.720 6.660 ;
        RECT 87.100 6.400 87.360 6.660 ;
        RECT 88.010 6.400 88.270 6.660 ;
        RECT 91.210 6.400 91.470 6.660 ;
        RECT 92.850 6.400 93.110 6.660 ;
        RECT 93.760 6.400 94.020 6.660 ;
        RECT 2.990 5.670 3.250 5.930 ;
        RECT 3.900 5.670 4.160 5.930 ;
        RECT 5.540 5.580 5.800 5.840 ;
        RECT 8.740 5.670 9.000 5.930 ;
        RECT 9.650 5.670 9.910 5.930 ;
        RECT 11.290 5.580 11.550 5.840 ;
        RECT 14.490 5.670 14.750 5.930 ;
        RECT 15.400 5.670 15.660 5.930 ;
        RECT 17.040 5.580 17.300 5.840 ;
        RECT 20.240 5.670 20.500 5.930 ;
        RECT 21.150 5.670 21.410 5.930 ;
        RECT 22.790 5.580 23.050 5.840 ;
        RECT 25.990 5.670 26.250 5.930 ;
        RECT 26.900 5.670 27.160 5.930 ;
        RECT 28.540 5.580 28.800 5.840 ;
        RECT 31.740 5.670 32.000 5.930 ;
        RECT 32.650 5.670 32.910 5.930 ;
        RECT 34.290 5.580 34.550 5.840 ;
        RECT 37.490 5.670 37.750 5.930 ;
        RECT 38.400 5.670 38.660 5.930 ;
        RECT 40.040 5.580 40.300 5.840 ;
        RECT 43.240 5.670 43.500 5.930 ;
        RECT 44.150 5.670 44.410 5.930 ;
        RECT 45.790 5.580 46.050 5.840 ;
        RECT 48.990 5.670 49.250 5.930 ;
        RECT 49.900 5.670 50.160 5.930 ;
        RECT 51.540 5.580 51.800 5.840 ;
        RECT 54.740 5.670 55.000 5.930 ;
        RECT 55.650 5.670 55.910 5.930 ;
        RECT 57.290 5.580 57.550 5.840 ;
        RECT 60.490 5.670 60.750 5.930 ;
        RECT 61.400 5.670 61.660 5.930 ;
        RECT 63.040 5.580 63.300 5.840 ;
        RECT 66.240 5.670 66.500 5.930 ;
        RECT 67.150 5.670 67.410 5.930 ;
        RECT 68.790 5.580 69.050 5.840 ;
        RECT 71.990 5.670 72.250 5.930 ;
        RECT 72.900 5.670 73.160 5.930 ;
        RECT 74.540 5.580 74.800 5.840 ;
        RECT 77.740 5.670 78.000 5.930 ;
        RECT 78.650 5.670 78.910 5.930 ;
        RECT 80.290 5.580 80.550 5.840 ;
        RECT 83.490 5.670 83.750 5.930 ;
        RECT 84.400 5.670 84.660 5.930 ;
        RECT 86.040 5.580 86.300 5.840 ;
        RECT 89.240 5.670 89.500 5.930 ;
        RECT 90.150 5.670 90.410 5.930 ;
        RECT 91.790 5.580 92.050 5.840 ;
        RECT 1.300 3.630 1.560 3.890 ;
        RECT 4.960 3.990 5.220 4.250 ;
        RECT 6.600 3.990 6.860 4.250 ;
        RECT 7.510 3.990 7.770 4.250 ;
        RECT 10.710 3.990 10.970 4.250 ;
        RECT 12.350 3.990 12.610 4.250 ;
        RECT 13.260 3.990 13.520 4.250 ;
        RECT 16.460 3.990 16.720 4.250 ;
        RECT 18.100 3.990 18.360 4.250 ;
        RECT 19.010 3.990 19.270 4.250 ;
        RECT 22.210 3.990 22.470 4.250 ;
        RECT 23.850 3.990 24.110 4.250 ;
        RECT 24.760 3.990 25.020 4.250 ;
        RECT 27.960 3.990 28.220 4.250 ;
        RECT 29.600 3.990 29.860 4.250 ;
        RECT 30.510 3.990 30.770 4.250 ;
        RECT 33.710 3.990 33.970 4.250 ;
        RECT 35.350 3.990 35.610 4.250 ;
        RECT 36.260 3.990 36.520 4.250 ;
        RECT 39.460 3.990 39.720 4.250 ;
        RECT 41.100 3.990 41.360 4.250 ;
        RECT 42.010 3.990 42.270 4.250 ;
        RECT 45.210 3.990 45.470 4.250 ;
        RECT 46.850 3.990 47.110 4.250 ;
        RECT 47.760 3.990 48.020 4.250 ;
        RECT 50.960 3.990 51.220 4.250 ;
        RECT 52.600 3.990 52.860 4.250 ;
        RECT 53.510 3.990 53.770 4.250 ;
        RECT 56.710 3.990 56.970 4.250 ;
        RECT 58.350 3.990 58.610 4.250 ;
        RECT 59.260 3.990 59.520 4.250 ;
        RECT 62.460 3.990 62.720 4.250 ;
        RECT 64.100 3.990 64.360 4.250 ;
        RECT 65.010 3.990 65.270 4.250 ;
        RECT 68.210 3.990 68.470 4.250 ;
        RECT 69.850 3.990 70.110 4.250 ;
        RECT 70.760 3.990 71.020 4.250 ;
        RECT 73.960 3.990 74.220 4.250 ;
        RECT 75.600 3.990 75.860 4.250 ;
        RECT 76.510 3.990 76.770 4.250 ;
        RECT 79.710 3.990 79.970 4.250 ;
        RECT 81.350 3.990 81.610 4.250 ;
        RECT 82.260 3.990 82.520 4.250 ;
        RECT 85.460 3.990 85.720 4.250 ;
        RECT 87.100 3.990 87.360 4.250 ;
        RECT 88.010 3.990 88.270 4.250 ;
        RECT 91.210 3.990 91.470 4.250 ;
        RECT 92.850 3.990 93.110 4.250 ;
        RECT 93.760 3.990 94.020 4.250 ;
        RECT 2.990 3.260 3.250 3.520 ;
        RECT 3.900 3.260 4.160 3.520 ;
        RECT 5.540 3.170 5.800 3.430 ;
        RECT 8.740 3.260 9.000 3.520 ;
        RECT 9.650 3.260 9.910 3.520 ;
        RECT 11.290 3.170 11.550 3.430 ;
        RECT 14.490 3.260 14.750 3.520 ;
        RECT 15.400 3.260 15.660 3.520 ;
        RECT 17.040 3.170 17.300 3.430 ;
        RECT 20.240 3.260 20.500 3.520 ;
        RECT 21.150 3.260 21.410 3.520 ;
        RECT 22.790 3.170 23.050 3.430 ;
        RECT 25.990 3.260 26.250 3.520 ;
        RECT 26.900 3.260 27.160 3.520 ;
        RECT 28.540 3.170 28.800 3.430 ;
        RECT 31.740 3.260 32.000 3.520 ;
        RECT 32.650 3.260 32.910 3.520 ;
        RECT 34.290 3.170 34.550 3.430 ;
        RECT 37.490 3.260 37.750 3.520 ;
        RECT 38.400 3.260 38.660 3.520 ;
        RECT 40.040 3.170 40.300 3.430 ;
        RECT 43.240 3.260 43.500 3.520 ;
        RECT 44.150 3.260 44.410 3.520 ;
        RECT 45.790 3.170 46.050 3.430 ;
        RECT 48.990 3.260 49.250 3.520 ;
        RECT 49.900 3.260 50.160 3.520 ;
        RECT 51.540 3.170 51.800 3.430 ;
        RECT 54.740 3.260 55.000 3.520 ;
        RECT 55.650 3.260 55.910 3.520 ;
        RECT 57.290 3.170 57.550 3.430 ;
        RECT 60.490 3.260 60.750 3.520 ;
        RECT 61.400 3.260 61.660 3.520 ;
        RECT 63.040 3.170 63.300 3.430 ;
        RECT 66.240 3.260 66.500 3.520 ;
        RECT 67.150 3.260 67.410 3.520 ;
        RECT 68.790 3.170 69.050 3.430 ;
        RECT 71.990 3.260 72.250 3.520 ;
        RECT 72.900 3.260 73.160 3.520 ;
        RECT 74.540 3.170 74.800 3.430 ;
        RECT 77.740 3.260 78.000 3.520 ;
        RECT 78.650 3.260 78.910 3.520 ;
        RECT 80.290 3.170 80.550 3.430 ;
        RECT 83.490 3.260 83.750 3.520 ;
        RECT 84.400 3.260 84.660 3.520 ;
        RECT 86.040 3.170 86.300 3.430 ;
        RECT 89.240 3.260 89.500 3.520 ;
        RECT 90.150 3.260 90.410 3.520 ;
        RECT 91.790 3.170 92.050 3.430 ;
        RECT 1.290 1.220 1.550 1.480 ;
        RECT 4.960 1.580 5.220 1.840 ;
        RECT 6.600 1.580 6.860 1.840 ;
        RECT 7.510 1.580 7.770 1.840 ;
        RECT 10.710 1.580 10.970 1.840 ;
        RECT 12.350 1.580 12.610 1.840 ;
        RECT 13.260 1.580 13.520 1.840 ;
        RECT 16.460 1.580 16.720 1.840 ;
        RECT 18.100 1.580 18.360 1.840 ;
        RECT 19.010 1.580 19.270 1.840 ;
        RECT 22.210 1.580 22.470 1.840 ;
        RECT 23.850 1.580 24.110 1.840 ;
        RECT 24.760 1.580 25.020 1.840 ;
        RECT 27.960 1.580 28.220 1.840 ;
        RECT 29.600 1.580 29.860 1.840 ;
        RECT 30.510 1.580 30.770 1.840 ;
        RECT 33.710 1.580 33.970 1.840 ;
        RECT 35.350 1.580 35.610 1.840 ;
        RECT 36.260 1.580 36.520 1.840 ;
        RECT 39.460 1.580 39.720 1.840 ;
        RECT 41.100 1.580 41.360 1.840 ;
        RECT 42.010 1.580 42.270 1.840 ;
        RECT 45.210 1.580 45.470 1.840 ;
        RECT 46.850 1.580 47.110 1.840 ;
        RECT 47.760 1.580 48.020 1.840 ;
        RECT 50.960 1.580 51.220 1.840 ;
        RECT 52.600 1.580 52.860 1.840 ;
        RECT 53.510 1.580 53.770 1.840 ;
        RECT 56.710 1.580 56.970 1.840 ;
        RECT 58.350 1.580 58.610 1.840 ;
        RECT 59.260 1.580 59.520 1.840 ;
        RECT 62.460 1.580 62.720 1.840 ;
        RECT 64.100 1.580 64.360 1.840 ;
        RECT 65.010 1.580 65.270 1.840 ;
        RECT 68.210 1.580 68.470 1.840 ;
        RECT 69.850 1.580 70.110 1.840 ;
        RECT 70.760 1.580 71.020 1.840 ;
        RECT 73.960 1.580 74.220 1.840 ;
        RECT 75.600 1.580 75.860 1.840 ;
        RECT 76.510 1.580 76.770 1.840 ;
        RECT 79.710 1.580 79.970 1.840 ;
        RECT 81.350 1.580 81.610 1.840 ;
        RECT 82.260 1.580 82.520 1.840 ;
        RECT 85.460 1.580 85.720 1.840 ;
        RECT 87.100 1.580 87.360 1.840 ;
        RECT 88.010 1.580 88.270 1.840 ;
        RECT 91.210 1.580 91.470 1.840 ;
        RECT 92.850 1.580 93.110 1.840 ;
        RECT 93.760 1.580 94.020 1.840 ;
        RECT 2.990 0.850 3.250 1.110 ;
        RECT 3.900 0.850 4.160 1.110 ;
        RECT 5.540 0.760 5.800 1.020 ;
        RECT 8.740 0.850 9.000 1.110 ;
        RECT 9.650 0.850 9.910 1.110 ;
        RECT 11.290 0.760 11.550 1.020 ;
        RECT 14.490 0.850 14.750 1.110 ;
        RECT 15.400 0.850 15.660 1.110 ;
        RECT 17.040 0.760 17.300 1.020 ;
        RECT 20.240 0.850 20.500 1.110 ;
        RECT 21.150 0.850 21.410 1.110 ;
        RECT 22.790 0.760 23.050 1.020 ;
        RECT 25.990 0.850 26.250 1.110 ;
        RECT 26.900 0.850 27.160 1.110 ;
        RECT 28.540 0.760 28.800 1.020 ;
        RECT 31.740 0.850 32.000 1.110 ;
        RECT 32.650 0.850 32.910 1.110 ;
        RECT 34.290 0.760 34.550 1.020 ;
        RECT 37.490 0.850 37.750 1.110 ;
        RECT 38.400 0.850 38.660 1.110 ;
        RECT 40.040 0.760 40.300 1.020 ;
        RECT 43.240 0.850 43.500 1.110 ;
        RECT 44.150 0.850 44.410 1.110 ;
        RECT 45.790 0.760 46.050 1.020 ;
        RECT 48.990 0.850 49.250 1.110 ;
        RECT 49.900 0.850 50.160 1.110 ;
        RECT 51.540 0.760 51.800 1.020 ;
        RECT 54.740 0.850 55.000 1.110 ;
        RECT 55.650 0.850 55.910 1.110 ;
        RECT 57.290 0.760 57.550 1.020 ;
        RECT 60.490 0.850 60.750 1.110 ;
        RECT 61.400 0.850 61.660 1.110 ;
        RECT 63.040 0.760 63.300 1.020 ;
        RECT 66.240 0.850 66.500 1.110 ;
        RECT 67.150 0.850 67.410 1.110 ;
        RECT 68.790 0.760 69.050 1.020 ;
        RECT 71.990 0.850 72.250 1.110 ;
        RECT 72.900 0.850 73.160 1.110 ;
        RECT 74.540 0.760 74.800 1.020 ;
        RECT 77.740 0.850 78.000 1.110 ;
        RECT 78.650 0.850 78.910 1.110 ;
        RECT 80.290 0.760 80.550 1.020 ;
        RECT 83.490 0.850 83.750 1.110 ;
        RECT 84.400 0.850 84.660 1.110 ;
        RECT 86.040 0.760 86.300 1.020 ;
        RECT 89.240 0.850 89.500 1.110 ;
        RECT 90.150 0.850 90.410 1.110 ;
        RECT 91.790 0.760 92.050 1.020 ;
        RECT 1.290 -1.190 1.550 -0.930 ;
        RECT 4.960 -0.830 5.220 -0.570 ;
        RECT 6.600 -0.830 6.860 -0.570 ;
        RECT 7.510 -0.830 7.770 -0.570 ;
        RECT 10.710 -0.830 10.970 -0.570 ;
        RECT 12.350 -0.830 12.610 -0.570 ;
        RECT 13.260 -0.830 13.520 -0.570 ;
        RECT 16.460 -0.830 16.720 -0.570 ;
        RECT 18.100 -0.830 18.360 -0.570 ;
        RECT 19.010 -0.830 19.270 -0.570 ;
        RECT 22.210 -0.830 22.470 -0.570 ;
        RECT 23.850 -0.830 24.110 -0.570 ;
        RECT 24.760 -0.830 25.020 -0.570 ;
        RECT 27.960 -0.830 28.220 -0.570 ;
        RECT 29.600 -0.830 29.860 -0.570 ;
        RECT 30.510 -0.830 30.770 -0.570 ;
        RECT 33.710 -0.830 33.970 -0.570 ;
        RECT 35.350 -0.830 35.610 -0.570 ;
        RECT 36.260 -0.830 36.520 -0.570 ;
        RECT 39.460 -0.830 39.720 -0.570 ;
        RECT 41.100 -0.830 41.360 -0.570 ;
        RECT 42.010 -0.830 42.270 -0.570 ;
        RECT 45.210 -0.830 45.470 -0.570 ;
        RECT 46.850 -0.830 47.110 -0.570 ;
        RECT 47.760 -0.830 48.020 -0.570 ;
        RECT 50.960 -0.830 51.220 -0.570 ;
        RECT 52.600 -0.830 52.860 -0.570 ;
        RECT 53.510 -0.830 53.770 -0.570 ;
        RECT 56.710 -0.830 56.970 -0.570 ;
        RECT 58.350 -0.830 58.610 -0.570 ;
        RECT 59.260 -0.830 59.520 -0.570 ;
        RECT 62.460 -0.830 62.720 -0.570 ;
        RECT 64.100 -0.830 64.360 -0.570 ;
        RECT 65.010 -0.830 65.270 -0.570 ;
        RECT 68.210 -0.830 68.470 -0.570 ;
        RECT 69.850 -0.830 70.110 -0.570 ;
        RECT 70.760 -0.830 71.020 -0.570 ;
        RECT 73.960 -0.830 74.220 -0.570 ;
        RECT 75.600 -0.830 75.860 -0.570 ;
        RECT 76.510 -0.830 76.770 -0.570 ;
        RECT 79.710 -0.830 79.970 -0.570 ;
        RECT 81.350 -0.830 81.610 -0.570 ;
        RECT 82.260 -0.830 82.520 -0.570 ;
        RECT 85.460 -0.830 85.720 -0.570 ;
        RECT 87.100 -0.830 87.360 -0.570 ;
        RECT 88.010 -0.830 88.270 -0.570 ;
        RECT 91.210 -0.830 91.470 -0.570 ;
        RECT 92.850 -0.830 93.110 -0.570 ;
        RECT 93.760 -0.830 94.020 -0.570 ;
        RECT 2.990 -1.560 3.250 -1.300 ;
        RECT 3.900 -1.560 4.160 -1.300 ;
        RECT 5.540 -1.650 5.800 -1.390 ;
        RECT 8.740 -1.560 9.000 -1.300 ;
        RECT 9.650 -1.560 9.910 -1.300 ;
        RECT 11.290 -1.650 11.550 -1.390 ;
        RECT 14.490 -1.560 14.750 -1.300 ;
        RECT 15.400 -1.560 15.660 -1.300 ;
        RECT 17.040 -1.650 17.300 -1.390 ;
        RECT 20.240 -1.560 20.500 -1.300 ;
        RECT 21.150 -1.560 21.410 -1.300 ;
        RECT 22.790 -1.650 23.050 -1.390 ;
        RECT 25.990 -1.560 26.250 -1.300 ;
        RECT 26.900 -1.560 27.160 -1.300 ;
        RECT 28.540 -1.650 28.800 -1.390 ;
        RECT 31.740 -1.560 32.000 -1.300 ;
        RECT 32.650 -1.560 32.910 -1.300 ;
        RECT 34.290 -1.650 34.550 -1.390 ;
        RECT 37.490 -1.560 37.750 -1.300 ;
        RECT 38.400 -1.560 38.660 -1.300 ;
        RECT 40.040 -1.650 40.300 -1.390 ;
        RECT 43.240 -1.560 43.500 -1.300 ;
        RECT 44.150 -1.560 44.410 -1.300 ;
        RECT 45.790 -1.650 46.050 -1.390 ;
        RECT 48.990 -1.560 49.250 -1.300 ;
        RECT 49.900 -1.560 50.160 -1.300 ;
        RECT 51.540 -1.650 51.800 -1.390 ;
        RECT 54.740 -1.560 55.000 -1.300 ;
        RECT 55.650 -1.560 55.910 -1.300 ;
        RECT 57.290 -1.650 57.550 -1.390 ;
        RECT 60.490 -1.560 60.750 -1.300 ;
        RECT 61.400 -1.560 61.660 -1.300 ;
        RECT 63.040 -1.650 63.300 -1.390 ;
        RECT 66.240 -1.560 66.500 -1.300 ;
        RECT 67.150 -1.560 67.410 -1.300 ;
        RECT 68.790 -1.650 69.050 -1.390 ;
        RECT 71.990 -1.560 72.250 -1.300 ;
        RECT 72.900 -1.560 73.160 -1.300 ;
        RECT 74.540 -1.650 74.800 -1.390 ;
        RECT 77.740 -1.560 78.000 -1.300 ;
        RECT 78.650 -1.560 78.910 -1.300 ;
        RECT 80.290 -1.650 80.550 -1.390 ;
        RECT 83.490 -1.560 83.750 -1.300 ;
        RECT 84.400 -1.560 84.660 -1.300 ;
        RECT 86.040 -1.650 86.300 -1.390 ;
        RECT 89.240 -1.560 89.500 -1.300 ;
        RECT 90.150 -1.560 90.410 -1.300 ;
        RECT 91.790 -1.650 92.050 -1.390 ;
        RECT 1.290 -2.040 1.550 -1.780 ;
        RECT 1.290 -2.830 1.550 -2.570 ;
        RECT 1.290 -3.600 1.550 -3.340 ;
        RECT 4.960 -3.240 5.220 -2.980 ;
        RECT 6.600 -3.240 6.860 -2.980 ;
        RECT 7.510 -3.240 7.770 -2.980 ;
        RECT 10.710 -3.240 10.970 -2.980 ;
        RECT 12.350 -3.240 12.610 -2.980 ;
        RECT 13.260 -3.240 13.520 -2.980 ;
        RECT 16.460 -3.240 16.720 -2.980 ;
        RECT 18.100 -3.240 18.360 -2.980 ;
        RECT 19.010 -3.240 19.270 -2.980 ;
        RECT 22.210 -3.240 22.470 -2.980 ;
        RECT 23.850 -3.240 24.110 -2.980 ;
        RECT 24.760 -3.240 25.020 -2.980 ;
        RECT 27.960 -3.240 28.220 -2.980 ;
        RECT 29.600 -3.240 29.860 -2.980 ;
        RECT 30.510 -3.240 30.770 -2.980 ;
        RECT 33.710 -3.240 33.970 -2.980 ;
        RECT 35.350 -3.240 35.610 -2.980 ;
        RECT 36.260 -3.240 36.520 -2.980 ;
        RECT 39.460 -3.240 39.720 -2.980 ;
        RECT 41.100 -3.240 41.360 -2.980 ;
        RECT 42.010 -3.240 42.270 -2.980 ;
        RECT 45.210 -3.240 45.470 -2.980 ;
        RECT 46.850 -3.240 47.110 -2.980 ;
        RECT 47.760 -3.240 48.020 -2.980 ;
        RECT 50.960 -3.240 51.220 -2.980 ;
        RECT 52.600 -3.240 52.860 -2.980 ;
        RECT 53.510 -3.240 53.770 -2.980 ;
        RECT 56.710 -3.240 56.970 -2.980 ;
        RECT 58.350 -3.240 58.610 -2.980 ;
        RECT 59.260 -3.240 59.520 -2.980 ;
        RECT 62.460 -3.240 62.720 -2.980 ;
        RECT 64.100 -3.240 64.360 -2.980 ;
        RECT 65.010 -3.240 65.270 -2.980 ;
        RECT 68.210 -3.240 68.470 -2.980 ;
        RECT 69.850 -3.240 70.110 -2.980 ;
        RECT 70.760 -3.240 71.020 -2.980 ;
        RECT 73.960 -3.240 74.220 -2.980 ;
        RECT 75.600 -3.240 75.860 -2.980 ;
        RECT 76.510 -3.240 76.770 -2.980 ;
        RECT 79.710 -3.240 79.970 -2.980 ;
        RECT 81.350 -3.240 81.610 -2.980 ;
        RECT 82.260 -3.240 82.520 -2.980 ;
        RECT 85.460 -3.240 85.720 -2.980 ;
        RECT 87.100 -3.240 87.360 -2.980 ;
        RECT 88.010 -3.240 88.270 -2.980 ;
        RECT 91.210 -3.240 91.470 -2.980 ;
        RECT 92.850 -3.240 93.110 -2.980 ;
        RECT 93.760 -3.240 94.020 -2.980 ;
        RECT 2.990 -3.970 3.250 -3.710 ;
        RECT 3.900 -3.970 4.160 -3.710 ;
        RECT 5.540 -4.060 5.800 -3.800 ;
        RECT 8.740 -3.970 9.000 -3.710 ;
        RECT 9.650 -3.970 9.910 -3.710 ;
        RECT 11.290 -4.060 11.550 -3.800 ;
        RECT 14.490 -3.970 14.750 -3.710 ;
        RECT 15.400 -3.970 15.660 -3.710 ;
        RECT 17.040 -4.060 17.300 -3.800 ;
        RECT 20.240 -3.970 20.500 -3.710 ;
        RECT 21.150 -3.970 21.410 -3.710 ;
        RECT 22.790 -4.060 23.050 -3.800 ;
        RECT 25.990 -3.970 26.250 -3.710 ;
        RECT 26.900 -3.970 27.160 -3.710 ;
        RECT 28.540 -4.060 28.800 -3.800 ;
        RECT 31.740 -3.970 32.000 -3.710 ;
        RECT 32.650 -3.970 32.910 -3.710 ;
        RECT 34.290 -4.060 34.550 -3.800 ;
        RECT 37.490 -3.970 37.750 -3.710 ;
        RECT 38.400 -3.970 38.660 -3.710 ;
        RECT 40.040 -4.060 40.300 -3.800 ;
        RECT 43.240 -3.970 43.500 -3.710 ;
        RECT 44.150 -3.970 44.410 -3.710 ;
        RECT 45.790 -4.060 46.050 -3.800 ;
        RECT 48.990 -3.970 49.250 -3.710 ;
        RECT 49.900 -3.970 50.160 -3.710 ;
        RECT 51.540 -4.060 51.800 -3.800 ;
        RECT 54.740 -3.970 55.000 -3.710 ;
        RECT 55.650 -3.970 55.910 -3.710 ;
        RECT 57.290 -4.060 57.550 -3.800 ;
        RECT 60.490 -3.970 60.750 -3.710 ;
        RECT 61.400 -3.970 61.660 -3.710 ;
        RECT 63.040 -4.060 63.300 -3.800 ;
        RECT 66.240 -3.970 66.500 -3.710 ;
        RECT 67.150 -3.970 67.410 -3.710 ;
        RECT 68.790 -4.060 69.050 -3.800 ;
        RECT 71.990 -3.970 72.250 -3.710 ;
        RECT 72.900 -3.970 73.160 -3.710 ;
        RECT 74.540 -4.060 74.800 -3.800 ;
        RECT 77.740 -3.970 78.000 -3.710 ;
        RECT 78.650 -3.970 78.910 -3.710 ;
        RECT 80.290 -4.060 80.550 -3.800 ;
        RECT 83.490 -3.970 83.750 -3.710 ;
        RECT 84.400 -3.970 84.660 -3.710 ;
        RECT 86.040 -4.060 86.300 -3.800 ;
        RECT 89.240 -3.970 89.500 -3.710 ;
        RECT 90.150 -3.970 90.410 -3.710 ;
        RECT 91.790 -4.060 92.050 -3.800 ;
        RECT 1.290 -4.420 1.550 -4.160 ;
        RECT 1.300 -5.210 1.560 -4.950 ;
        RECT 1.290 -6.010 1.550 -5.750 ;
        RECT 4.960 -5.650 5.220 -5.390 ;
        RECT 6.600 -5.650 6.860 -5.390 ;
        RECT 7.510 -5.650 7.770 -5.390 ;
        RECT 10.710 -5.650 10.970 -5.390 ;
        RECT 12.350 -5.650 12.610 -5.390 ;
        RECT 13.260 -5.650 13.520 -5.390 ;
        RECT 16.460 -5.650 16.720 -5.390 ;
        RECT 18.100 -5.650 18.360 -5.390 ;
        RECT 19.010 -5.650 19.270 -5.390 ;
        RECT 22.210 -5.650 22.470 -5.390 ;
        RECT 23.850 -5.650 24.110 -5.390 ;
        RECT 24.760 -5.650 25.020 -5.390 ;
        RECT 27.960 -5.650 28.220 -5.390 ;
        RECT 29.600 -5.650 29.860 -5.390 ;
        RECT 30.510 -5.650 30.770 -5.390 ;
        RECT 33.710 -5.650 33.970 -5.390 ;
        RECT 35.350 -5.650 35.610 -5.390 ;
        RECT 36.260 -5.650 36.520 -5.390 ;
        RECT 39.460 -5.650 39.720 -5.390 ;
        RECT 41.100 -5.650 41.360 -5.390 ;
        RECT 42.010 -5.650 42.270 -5.390 ;
        RECT 45.210 -5.650 45.470 -5.390 ;
        RECT 46.850 -5.650 47.110 -5.390 ;
        RECT 47.760 -5.650 48.020 -5.390 ;
        RECT 50.960 -5.650 51.220 -5.390 ;
        RECT 52.600 -5.650 52.860 -5.390 ;
        RECT 53.510 -5.650 53.770 -5.390 ;
        RECT 56.710 -5.650 56.970 -5.390 ;
        RECT 58.350 -5.650 58.610 -5.390 ;
        RECT 59.260 -5.650 59.520 -5.390 ;
        RECT 62.460 -5.650 62.720 -5.390 ;
        RECT 64.100 -5.650 64.360 -5.390 ;
        RECT 65.010 -5.650 65.270 -5.390 ;
        RECT 68.210 -5.650 68.470 -5.390 ;
        RECT 69.850 -5.650 70.110 -5.390 ;
        RECT 70.760 -5.650 71.020 -5.390 ;
        RECT 73.960 -5.650 74.220 -5.390 ;
        RECT 75.600 -5.650 75.860 -5.390 ;
        RECT 76.510 -5.650 76.770 -5.390 ;
        RECT 79.710 -5.650 79.970 -5.390 ;
        RECT 81.350 -5.650 81.610 -5.390 ;
        RECT 82.260 -5.650 82.520 -5.390 ;
        RECT 85.460 -5.650 85.720 -5.390 ;
        RECT 87.100 -5.650 87.360 -5.390 ;
        RECT 88.010 -5.650 88.270 -5.390 ;
        RECT 91.210 -5.650 91.470 -5.390 ;
        RECT 92.850 -5.650 93.110 -5.390 ;
        RECT 93.760 -5.650 94.020 -5.390 ;
        RECT 2.990 -6.970 3.250 -6.710 ;
        RECT 3.900 -6.970 4.160 -6.710 ;
        RECT 5.540 -7.060 5.800 -6.800 ;
        RECT 8.740 -6.970 9.000 -6.710 ;
        RECT 9.650 -6.970 9.910 -6.710 ;
        RECT 11.290 -7.060 11.550 -6.800 ;
        RECT 14.490 -6.970 14.750 -6.710 ;
        RECT 15.400 -6.970 15.660 -6.710 ;
        RECT 17.040 -7.060 17.300 -6.800 ;
        RECT 20.240 -6.970 20.500 -6.710 ;
        RECT 21.150 -6.970 21.410 -6.710 ;
        RECT 22.790 -7.060 23.050 -6.800 ;
        RECT 25.990 -6.970 26.250 -6.710 ;
        RECT 26.900 -6.970 27.160 -6.710 ;
        RECT 28.540 -7.060 28.800 -6.800 ;
        RECT 31.740 -6.970 32.000 -6.710 ;
        RECT 32.650 -6.970 32.910 -6.710 ;
        RECT 34.290 -7.060 34.550 -6.800 ;
        RECT 37.490 -6.970 37.750 -6.710 ;
        RECT 38.400 -6.970 38.660 -6.710 ;
        RECT 40.040 -7.060 40.300 -6.800 ;
        RECT 43.240 -6.970 43.500 -6.710 ;
        RECT 44.150 -6.970 44.410 -6.710 ;
        RECT 45.790 -7.060 46.050 -6.800 ;
        RECT 48.990 -6.970 49.250 -6.710 ;
        RECT 49.900 -6.970 50.160 -6.710 ;
        RECT 51.540 -7.060 51.800 -6.800 ;
        RECT 54.740 -6.970 55.000 -6.710 ;
        RECT 55.650 -6.970 55.910 -6.710 ;
        RECT 57.290 -7.060 57.550 -6.800 ;
        RECT 60.490 -6.970 60.750 -6.710 ;
        RECT 61.400 -6.970 61.660 -6.710 ;
        RECT 63.040 -7.060 63.300 -6.800 ;
        RECT 66.240 -6.970 66.500 -6.710 ;
        RECT 67.150 -6.970 67.410 -6.710 ;
        RECT 68.790 -7.060 69.050 -6.800 ;
        RECT 71.990 -6.970 72.250 -6.710 ;
        RECT 72.900 -6.970 73.160 -6.710 ;
        RECT 74.540 -7.060 74.800 -6.800 ;
        RECT 77.740 -6.970 78.000 -6.710 ;
        RECT 78.650 -6.970 78.910 -6.710 ;
        RECT 80.290 -7.060 80.550 -6.800 ;
        RECT 83.490 -6.970 83.750 -6.710 ;
        RECT 84.400 -6.970 84.660 -6.710 ;
        RECT 86.040 -7.060 86.300 -6.800 ;
        RECT 89.240 -6.970 89.500 -6.710 ;
        RECT 90.150 -6.970 90.410 -6.710 ;
        RECT 91.790 -7.060 92.050 -6.800 ;
        RECT 1.290 -7.440 1.550 -7.180 ;
        RECT 1.290 -8.240 1.550 -7.980 ;
        RECT 1.290 -9.010 1.550 -8.750 ;
        RECT 4.960 -8.650 5.220 -8.390 ;
        RECT 6.600 -8.650 6.860 -8.390 ;
        RECT 7.510 -8.650 7.770 -8.390 ;
        RECT 10.710 -8.650 10.970 -8.390 ;
        RECT 12.350 -8.650 12.610 -8.390 ;
        RECT 13.260 -8.650 13.520 -8.390 ;
        RECT 16.460 -8.650 16.720 -8.390 ;
        RECT 18.100 -8.650 18.360 -8.390 ;
        RECT 19.010 -8.650 19.270 -8.390 ;
        RECT 22.210 -8.650 22.470 -8.390 ;
        RECT 23.850 -8.650 24.110 -8.390 ;
        RECT 24.760 -8.650 25.020 -8.390 ;
        RECT 27.960 -8.650 28.220 -8.390 ;
        RECT 29.600 -8.650 29.860 -8.390 ;
        RECT 30.510 -8.650 30.770 -8.390 ;
        RECT 33.710 -8.650 33.970 -8.390 ;
        RECT 35.350 -8.650 35.610 -8.390 ;
        RECT 36.260 -8.650 36.520 -8.390 ;
        RECT 39.460 -8.650 39.720 -8.390 ;
        RECT 41.100 -8.650 41.360 -8.390 ;
        RECT 42.010 -8.650 42.270 -8.390 ;
        RECT 45.210 -8.650 45.470 -8.390 ;
        RECT 46.850 -8.650 47.110 -8.390 ;
        RECT 47.760 -8.650 48.020 -8.390 ;
        RECT 50.960 -8.650 51.220 -8.390 ;
        RECT 52.600 -8.650 52.860 -8.390 ;
        RECT 53.510 -8.650 53.770 -8.390 ;
        RECT 56.710 -8.650 56.970 -8.390 ;
        RECT 58.350 -8.650 58.610 -8.390 ;
        RECT 59.260 -8.650 59.520 -8.390 ;
        RECT 62.460 -8.650 62.720 -8.390 ;
        RECT 64.100 -8.650 64.360 -8.390 ;
        RECT 65.010 -8.650 65.270 -8.390 ;
        RECT 68.210 -8.650 68.470 -8.390 ;
        RECT 69.850 -8.650 70.110 -8.390 ;
        RECT 70.760 -8.650 71.020 -8.390 ;
        RECT 73.960 -8.650 74.220 -8.390 ;
        RECT 75.600 -8.650 75.860 -8.390 ;
        RECT 76.510 -8.650 76.770 -8.390 ;
        RECT 79.710 -8.650 79.970 -8.390 ;
        RECT 81.350 -8.650 81.610 -8.390 ;
        RECT 82.260 -8.650 82.520 -8.390 ;
        RECT 85.460 -8.650 85.720 -8.390 ;
        RECT 87.100 -8.650 87.360 -8.390 ;
        RECT 88.010 -8.650 88.270 -8.390 ;
        RECT 91.210 -8.650 91.470 -8.390 ;
        RECT 92.850 -8.650 93.110 -8.390 ;
        RECT 93.760 -8.650 94.020 -8.390 ;
        RECT 2.990 -9.380 3.250 -9.120 ;
        RECT 3.900 -9.380 4.160 -9.120 ;
        RECT 5.540 -9.470 5.800 -9.210 ;
        RECT 8.740 -9.380 9.000 -9.120 ;
        RECT 9.650 -9.380 9.910 -9.120 ;
        RECT 11.290 -9.470 11.550 -9.210 ;
        RECT 14.490 -9.380 14.750 -9.120 ;
        RECT 15.400 -9.380 15.660 -9.120 ;
        RECT 17.040 -9.470 17.300 -9.210 ;
        RECT 20.240 -9.380 20.500 -9.120 ;
        RECT 21.150 -9.380 21.410 -9.120 ;
        RECT 22.790 -9.470 23.050 -9.210 ;
        RECT 25.990 -9.380 26.250 -9.120 ;
        RECT 26.900 -9.380 27.160 -9.120 ;
        RECT 28.540 -9.470 28.800 -9.210 ;
        RECT 31.740 -9.380 32.000 -9.120 ;
        RECT 32.650 -9.380 32.910 -9.120 ;
        RECT 34.290 -9.470 34.550 -9.210 ;
        RECT 37.490 -9.380 37.750 -9.120 ;
        RECT 38.400 -9.380 38.660 -9.120 ;
        RECT 40.040 -9.470 40.300 -9.210 ;
        RECT 43.240 -9.380 43.500 -9.120 ;
        RECT 44.150 -9.380 44.410 -9.120 ;
        RECT 45.790 -9.470 46.050 -9.210 ;
        RECT 48.990 -9.380 49.250 -9.120 ;
        RECT 49.900 -9.380 50.160 -9.120 ;
        RECT 51.540 -9.470 51.800 -9.210 ;
        RECT 54.740 -9.380 55.000 -9.120 ;
        RECT 55.650 -9.380 55.910 -9.120 ;
        RECT 57.290 -9.470 57.550 -9.210 ;
        RECT 60.490 -9.380 60.750 -9.120 ;
        RECT 61.400 -9.380 61.660 -9.120 ;
        RECT 63.040 -9.470 63.300 -9.210 ;
        RECT 66.240 -9.380 66.500 -9.120 ;
        RECT 67.150 -9.380 67.410 -9.120 ;
        RECT 68.790 -9.470 69.050 -9.210 ;
        RECT 71.990 -9.380 72.250 -9.120 ;
        RECT 72.900 -9.380 73.160 -9.120 ;
        RECT 74.540 -9.470 74.800 -9.210 ;
        RECT 77.740 -9.380 78.000 -9.120 ;
        RECT 78.650 -9.380 78.910 -9.120 ;
        RECT 80.290 -9.470 80.550 -9.210 ;
        RECT 83.490 -9.380 83.750 -9.120 ;
        RECT 84.400 -9.380 84.660 -9.120 ;
        RECT 86.040 -9.470 86.300 -9.210 ;
        RECT 89.240 -9.380 89.500 -9.120 ;
        RECT 90.150 -9.380 90.410 -9.120 ;
        RECT 91.790 -9.470 92.050 -9.210 ;
        RECT 1.290 -9.810 1.550 -9.550 ;
        RECT 1.300 -10.680 1.560 -10.420 ;
        RECT 1.290 -11.420 1.550 -11.160 ;
        RECT 4.960 -11.060 5.220 -10.800 ;
        RECT 6.600 -11.060 6.860 -10.800 ;
        RECT 7.510 -11.060 7.770 -10.800 ;
        RECT 10.710 -11.060 10.970 -10.800 ;
        RECT 12.350 -11.060 12.610 -10.800 ;
        RECT 13.260 -11.060 13.520 -10.800 ;
        RECT 16.460 -11.060 16.720 -10.800 ;
        RECT 18.100 -11.060 18.360 -10.800 ;
        RECT 19.010 -11.060 19.270 -10.800 ;
        RECT 22.210 -11.060 22.470 -10.800 ;
        RECT 23.850 -11.060 24.110 -10.800 ;
        RECT 24.760 -11.060 25.020 -10.800 ;
        RECT 27.960 -11.060 28.220 -10.800 ;
        RECT 29.600 -11.060 29.860 -10.800 ;
        RECT 30.510 -11.060 30.770 -10.800 ;
        RECT 33.710 -11.060 33.970 -10.800 ;
        RECT 35.350 -11.060 35.610 -10.800 ;
        RECT 36.260 -11.060 36.520 -10.800 ;
        RECT 39.460 -11.060 39.720 -10.800 ;
        RECT 41.100 -11.060 41.360 -10.800 ;
        RECT 42.010 -11.060 42.270 -10.800 ;
        RECT 45.210 -11.060 45.470 -10.800 ;
        RECT 46.850 -11.060 47.110 -10.800 ;
        RECT 47.760 -11.060 48.020 -10.800 ;
        RECT 50.960 -11.060 51.220 -10.800 ;
        RECT 52.600 -11.060 52.860 -10.800 ;
        RECT 53.510 -11.060 53.770 -10.800 ;
        RECT 56.710 -11.060 56.970 -10.800 ;
        RECT 58.350 -11.060 58.610 -10.800 ;
        RECT 59.260 -11.060 59.520 -10.800 ;
        RECT 62.460 -11.060 62.720 -10.800 ;
        RECT 64.100 -11.060 64.360 -10.800 ;
        RECT 65.010 -11.060 65.270 -10.800 ;
        RECT 68.210 -11.060 68.470 -10.800 ;
        RECT 69.850 -11.060 70.110 -10.800 ;
        RECT 70.760 -11.060 71.020 -10.800 ;
        RECT 73.960 -11.060 74.220 -10.800 ;
        RECT 75.600 -11.060 75.860 -10.800 ;
        RECT 76.510 -11.060 76.770 -10.800 ;
        RECT 79.710 -11.060 79.970 -10.800 ;
        RECT 81.350 -11.060 81.610 -10.800 ;
        RECT 82.260 -11.060 82.520 -10.800 ;
        RECT 85.460 -11.060 85.720 -10.800 ;
        RECT 87.100 -11.060 87.360 -10.800 ;
        RECT 88.010 -11.060 88.270 -10.800 ;
        RECT 91.210 -11.060 91.470 -10.800 ;
        RECT 92.850 -11.060 93.110 -10.800 ;
        RECT 93.760 -11.060 94.020 -10.800 ;
        RECT 5.260 -12.880 5.520 -12.620 ;
        RECT 11.010 -12.880 11.270 -12.620 ;
        RECT 16.760 -12.880 17.020 -12.620 ;
        RECT 22.510 -12.880 22.770 -12.620 ;
        RECT 28.260 -12.880 28.520 -12.620 ;
        RECT 34.010 -12.880 34.270 -12.620 ;
        RECT 39.760 -12.880 40.020 -12.620 ;
        RECT 45.510 -12.880 45.770 -12.620 ;
        RECT 51.260 -12.880 51.520 -12.620 ;
        RECT 57.010 -12.880 57.270 -12.620 ;
        RECT 62.760 -12.880 63.020 -12.620 ;
        RECT 68.510 -12.880 68.770 -12.620 ;
        RECT 74.260 -12.880 74.520 -12.620 ;
        RECT 80.010 -12.880 80.270 -12.620 ;
        RECT 85.760 -12.880 86.020 -12.620 ;
        RECT 91.510 -12.880 91.770 -12.620 ;
        RECT 5.970 -14.120 6.230 -13.860 ;
        RECT 11.720 -14.130 11.980 -13.870 ;
        RECT 17.470 -14.150 17.730 -13.890 ;
        RECT 23.220 -14.150 23.480 -13.890 ;
        RECT 28.970 -14.130 29.230 -13.870 ;
        RECT 34.720 -14.100 34.980 -13.840 ;
        RECT 40.470 -14.080 40.730 -13.820 ;
        RECT 46.220 -14.080 46.480 -13.820 ;
        RECT 51.970 -14.130 52.230 -13.870 ;
        RECT 57.720 -14.100 57.980 -13.840 ;
        RECT 63.470 -14.140 63.730 -13.880 ;
        RECT 69.220 -14.150 69.480 -13.890 ;
        RECT 74.970 -14.110 75.230 -13.850 ;
        RECT 80.720 -14.150 80.980 -13.890 ;
        RECT 86.470 -14.110 86.730 -13.850 ;
        RECT 92.220 -14.120 92.480 -13.860 ;
        RECT 3.360 -14.540 3.620 -14.280 ;
        RECT 3.900 -14.540 4.160 -14.280 ;
        RECT 6.610 -14.540 6.870 -14.280 ;
        RECT 7.150 -14.540 7.410 -14.280 ;
        RECT 9.110 -14.540 9.370 -14.280 ;
        RECT 9.650 -14.540 9.910 -14.280 ;
        RECT 12.360 -14.540 12.620 -14.280 ;
        RECT 12.900 -14.540 13.160 -14.280 ;
        RECT 14.860 -14.540 15.120 -14.280 ;
        RECT 15.400 -14.540 15.660 -14.280 ;
        RECT 18.110 -14.540 18.370 -14.280 ;
        RECT 18.650 -14.540 18.910 -14.280 ;
        RECT 20.610 -14.540 20.870 -14.280 ;
        RECT 21.150 -14.540 21.410 -14.280 ;
        RECT 23.860 -14.540 24.120 -14.280 ;
        RECT 24.400 -14.540 24.660 -14.280 ;
        RECT 26.360 -14.540 26.620 -14.280 ;
        RECT 26.900 -14.540 27.160 -14.280 ;
        RECT 29.610 -14.540 29.870 -14.280 ;
        RECT 30.150 -14.540 30.410 -14.280 ;
        RECT 32.110 -14.540 32.370 -14.280 ;
        RECT 32.650 -14.540 32.910 -14.280 ;
        RECT 35.360 -14.540 35.620 -14.280 ;
        RECT 35.900 -14.540 36.160 -14.280 ;
        RECT 37.860 -14.540 38.120 -14.280 ;
        RECT 38.400 -14.540 38.660 -14.280 ;
        RECT 41.110 -14.540 41.370 -14.280 ;
        RECT 41.650 -14.540 41.910 -14.280 ;
        RECT 43.610 -14.540 43.870 -14.280 ;
        RECT 44.150 -14.540 44.410 -14.280 ;
        RECT 46.860 -14.540 47.120 -14.280 ;
        RECT 47.400 -14.540 47.660 -14.280 ;
        RECT 49.360 -14.540 49.620 -14.280 ;
        RECT 49.900 -14.540 50.160 -14.280 ;
        RECT 52.610 -14.540 52.870 -14.280 ;
        RECT 53.150 -14.540 53.410 -14.280 ;
        RECT 55.110 -14.540 55.370 -14.280 ;
        RECT 55.650 -14.540 55.910 -14.280 ;
        RECT 58.360 -14.540 58.620 -14.280 ;
        RECT 58.900 -14.540 59.160 -14.280 ;
        RECT 60.860 -14.540 61.120 -14.280 ;
        RECT 61.400 -14.540 61.660 -14.280 ;
        RECT 64.110 -14.540 64.370 -14.280 ;
        RECT 64.650 -14.540 64.910 -14.280 ;
        RECT 66.610 -14.540 66.870 -14.280 ;
        RECT 67.150 -14.540 67.410 -14.280 ;
        RECT 69.860 -14.540 70.120 -14.280 ;
        RECT 70.400 -14.540 70.660 -14.280 ;
        RECT 72.360 -14.540 72.620 -14.280 ;
        RECT 72.900 -14.540 73.160 -14.280 ;
        RECT 75.610 -14.540 75.870 -14.280 ;
        RECT 76.150 -14.540 76.410 -14.280 ;
        RECT 78.110 -14.540 78.370 -14.280 ;
        RECT 78.650 -14.540 78.910 -14.280 ;
        RECT 81.360 -14.540 81.620 -14.280 ;
        RECT 81.900 -14.540 82.160 -14.280 ;
        RECT 83.860 -14.540 84.120 -14.280 ;
        RECT 84.400 -14.540 84.660 -14.280 ;
        RECT 87.110 -14.540 87.370 -14.280 ;
        RECT 87.650 -14.540 87.910 -14.280 ;
        RECT 89.610 -14.540 89.870 -14.280 ;
        RECT 90.150 -14.540 90.410 -14.280 ;
        RECT 92.860 -14.540 93.120 -14.280 ;
        RECT 93.400 -14.540 93.660 -14.280 ;
        RECT 3.430 -18.740 3.690 -18.480 ;
        RECT 7.110 -18.750 7.370 -18.490 ;
        RECT 9.180 -18.740 9.440 -18.480 ;
        RECT 12.860 -18.750 13.120 -18.490 ;
        RECT 14.930 -18.740 15.190 -18.480 ;
        RECT 18.610 -18.750 18.870 -18.490 ;
        RECT 20.680 -18.740 20.940 -18.480 ;
        RECT 24.360 -18.750 24.620 -18.490 ;
        RECT 26.430 -18.740 26.690 -18.480 ;
        RECT 30.110 -18.750 30.370 -18.490 ;
        RECT 32.180 -18.740 32.440 -18.480 ;
        RECT 35.860 -18.750 36.120 -18.490 ;
        RECT 37.930 -18.740 38.190 -18.480 ;
        RECT 41.610 -18.750 41.870 -18.490 ;
        RECT 43.680 -18.740 43.940 -18.480 ;
        RECT 47.360 -18.750 47.620 -18.490 ;
        RECT 49.430 -18.740 49.690 -18.480 ;
        RECT 53.110 -18.750 53.370 -18.490 ;
        RECT 55.180 -18.740 55.440 -18.480 ;
        RECT 58.860 -18.750 59.120 -18.490 ;
        RECT 60.930 -18.740 61.190 -18.480 ;
        RECT 64.610 -18.750 64.870 -18.490 ;
        RECT 66.680 -18.740 66.940 -18.480 ;
        RECT 70.360 -18.750 70.620 -18.490 ;
        RECT 72.430 -18.740 72.690 -18.480 ;
        RECT 76.110 -18.750 76.370 -18.490 ;
        RECT 78.180 -18.740 78.440 -18.480 ;
        RECT 81.860 -18.750 82.120 -18.490 ;
        RECT 83.930 -18.740 84.190 -18.480 ;
        RECT 87.610 -18.750 87.870 -18.490 ;
        RECT 89.680 -18.740 89.940 -18.480 ;
        RECT 93.360 -18.750 93.620 -18.490 ;
        RECT 1.290 -19.190 1.550 -18.930 ;
        RECT 4.110 -20.180 4.370 -19.920 ;
        RECT 6.390 -20.180 6.650 -19.920 ;
        RECT 9.860 -20.180 10.120 -19.920 ;
        RECT 12.140 -20.180 12.400 -19.920 ;
        RECT 15.610 -20.180 15.870 -19.920 ;
        RECT 17.890 -20.180 18.150 -19.920 ;
        RECT 21.360 -20.180 21.620 -19.920 ;
        RECT 23.640 -20.180 23.900 -19.920 ;
        RECT 27.110 -20.180 27.370 -19.920 ;
        RECT 29.390 -20.180 29.650 -19.920 ;
        RECT 32.860 -20.180 33.120 -19.920 ;
        RECT 35.140 -20.180 35.400 -19.920 ;
        RECT 38.610 -20.180 38.870 -19.920 ;
        RECT 40.890 -20.180 41.150 -19.920 ;
        RECT 44.360 -20.180 44.620 -19.920 ;
        RECT 46.640 -20.180 46.900 -19.920 ;
        RECT 50.110 -20.180 50.370 -19.920 ;
        RECT 52.390 -20.180 52.650 -19.920 ;
        RECT 55.860 -20.180 56.120 -19.920 ;
        RECT 58.140 -20.180 58.400 -19.920 ;
        RECT 61.610 -20.180 61.870 -19.920 ;
        RECT 63.890 -20.180 64.150 -19.920 ;
        RECT 67.360 -20.180 67.620 -19.920 ;
        RECT 69.640 -20.180 69.900 -19.920 ;
        RECT 73.110 -20.180 73.370 -19.920 ;
        RECT 75.390 -20.180 75.650 -19.920 ;
        RECT 78.860 -20.180 79.120 -19.920 ;
        RECT 81.140 -20.180 81.400 -19.920 ;
        RECT 84.610 -20.180 84.870 -19.920 ;
        RECT 86.890 -20.180 87.150 -19.920 ;
        RECT 90.360 -20.180 90.620 -19.920 ;
        RECT 92.640 -20.180 92.900 -19.920 ;
        RECT -0.330 -20.580 -0.070 -20.320 ;
        RECT 1.300 -20.590 1.560 -20.330 ;
        RECT 2.280 -21.270 2.540 -21.010 ;
        RECT 8.090 -21.250 8.350 -20.990 ;
        RECT 13.810 -21.260 14.070 -21.000 ;
        RECT 19.590 -21.280 19.850 -21.020 ;
        RECT 25.340 -21.280 25.600 -21.020 ;
        RECT 31.050 -21.300 31.310 -21.040 ;
        RECT 36.820 -21.290 37.080 -21.030 ;
        RECT 42.620 -21.280 42.880 -21.020 ;
        RECT 48.320 -21.270 48.580 -21.010 ;
        RECT 54.090 -21.290 54.350 -21.030 ;
        RECT 59.830 -21.270 60.090 -21.010 ;
        RECT 65.560 -21.280 65.820 -21.020 ;
        RECT 71.330 -21.290 71.590 -21.030 ;
        RECT 77.090 -21.290 77.350 -21.030 ;
        RECT 82.820 -21.310 83.080 -21.050 ;
        RECT 88.570 -21.310 88.830 -21.050 ;
        RECT 5.260 -22.070 5.520 -21.810 ;
        RECT 11.010 -22.070 11.270 -21.810 ;
        RECT 16.760 -22.070 17.020 -21.810 ;
        RECT 22.510 -22.070 22.770 -21.810 ;
        RECT 28.260 -22.070 28.520 -21.810 ;
        RECT 34.010 -22.070 34.270 -21.810 ;
        RECT 39.760 -22.070 40.020 -21.810 ;
        RECT 45.510 -22.070 45.770 -21.810 ;
        RECT 51.260 -22.070 51.520 -21.810 ;
        RECT 57.010 -22.070 57.270 -21.810 ;
        RECT 62.760 -22.070 63.020 -21.810 ;
        RECT 68.510 -22.070 68.770 -21.810 ;
        RECT 74.260 -22.070 74.520 -21.810 ;
        RECT 80.010 -22.070 80.270 -21.810 ;
        RECT 85.760 -22.070 86.020 -21.810 ;
        RECT 91.510 -22.070 91.770 -21.810 ;
        RECT 2.990 -23.000 3.250 -22.740 ;
        RECT 7.520 -23.000 7.780 -22.740 ;
        RECT 8.740 -23.000 9.000 -22.740 ;
        RECT 13.270 -23.000 13.530 -22.740 ;
        RECT 14.490 -23.000 14.750 -22.740 ;
        RECT 19.020 -23.000 19.280 -22.740 ;
        RECT 20.240 -23.000 20.500 -22.740 ;
        RECT 24.770 -23.000 25.030 -22.740 ;
        RECT 25.990 -23.000 26.250 -22.740 ;
        RECT 30.520 -23.000 30.780 -22.740 ;
        RECT 31.740 -23.000 32.000 -22.740 ;
        RECT 36.270 -23.000 36.530 -22.740 ;
        RECT 37.490 -23.000 37.750 -22.740 ;
        RECT 42.020 -23.000 42.280 -22.740 ;
        RECT 43.240 -23.000 43.500 -22.740 ;
        RECT 47.770 -23.000 48.030 -22.740 ;
        RECT 48.990 -23.000 49.250 -22.740 ;
        RECT 53.520 -23.000 53.780 -22.740 ;
        RECT 54.740 -23.000 55.000 -22.740 ;
        RECT 59.270 -23.000 59.530 -22.740 ;
        RECT 60.490 -23.000 60.750 -22.740 ;
        RECT 65.020 -23.000 65.280 -22.740 ;
        RECT 66.240 -23.000 66.500 -22.740 ;
        RECT 70.770 -23.000 71.030 -22.740 ;
        RECT 71.990 -23.000 72.250 -22.740 ;
        RECT 76.520 -23.000 76.780 -22.740 ;
        RECT 77.740 -23.000 78.000 -22.740 ;
        RECT 82.270 -23.000 82.530 -22.740 ;
        RECT 83.490 -23.000 83.750 -22.740 ;
        RECT 88.020 -23.000 88.280 -22.740 ;
        RECT 89.240 -23.000 89.500 -22.740 ;
        RECT 93.770 -23.000 94.030 -22.740 ;
        RECT 5.260 -23.670 5.520 -23.410 ;
        RECT 8.130 -23.480 8.390 -23.220 ;
        RECT 11.010 -23.680 11.270 -23.420 ;
        RECT 16.760 -23.730 17.020 -23.470 ;
        RECT 19.620 -23.490 19.880 -23.230 ;
        RECT 22.510 -23.730 22.770 -23.470 ;
        RECT 28.260 -23.730 28.520 -23.470 ;
        RECT 31.050 -23.500 31.310 -23.240 ;
        RECT 34.010 -23.730 34.270 -23.470 ;
        RECT 39.760 -23.730 40.020 -23.470 ;
        RECT 42.620 -23.510 42.880 -23.250 ;
        RECT 45.510 -23.730 45.770 -23.470 ;
        RECT 51.260 -23.730 51.520 -23.470 ;
        RECT 54.020 -23.490 54.280 -23.230 ;
        RECT 57.010 -23.730 57.270 -23.470 ;
        RECT 62.760 -23.730 63.020 -23.470 ;
        RECT 65.700 -23.490 65.960 -23.230 ;
        RECT 68.510 -23.730 68.770 -23.470 ;
        RECT 74.260 -23.730 74.520 -23.470 ;
        RECT 77.150 -23.490 77.410 -23.230 ;
        RECT 88.720 -23.470 88.980 -23.210 ;
        RECT 80.010 -23.730 80.270 -23.470 ;
        RECT 85.760 -23.730 86.020 -23.470 ;
        RECT 91.510 -23.730 91.770 -23.470 ;
        RECT 7.370 -24.470 7.630 -24.210 ;
        RECT 8.920 -24.470 9.180 -24.210 ;
        RECT 18.870 -24.470 19.130 -24.210 ;
        RECT 20.420 -24.470 20.680 -24.210 ;
        RECT 30.370 -24.470 30.630 -24.210 ;
        RECT 31.910 -24.470 32.170 -24.210 ;
        RECT 41.840 -24.470 42.100 -24.210 ;
        RECT 43.430 -24.480 43.690 -24.220 ;
        RECT -39.240 -24.840 -38.980 -24.580 ;
        RECT 53.360 -24.470 53.620 -24.210 ;
        RECT 54.910 -24.470 55.170 -24.210 ;
        RECT 64.870 -24.480 65.130 -24.220 ;
        RECT 66.400 -24.480 66.660 -24.220 ;
        RECT 76.380 -24.470 76.640 -24.210 ;
        RECT 77.910 -24.470 78.170 -24.210 ;
        RECT 87.870 -24.460 88.130 -24.200 ;
        RECT 89.390 -24.470 89.650 -24.210 ;
        RECT 4.680 -25.240 4.940 -24.980 ;
        RECT 11.610 -25.170 11.870 -24.910 ;
        RECT 16.170 -25.160 16.430 -24.900 ;
        RECT 23.100 -25.210 23.360 -24.950 ;
        RECT 27.690 -25.220 27.950 -24.960 ;
        RECT 34.610 -25.200 34.870 -24.940 ;
        RECT 39.190 -25.220 39.450 -24.960 ;
        RECT 46.100 -25.240 46.360 -24.980 ;
        RECT 50.680 -25.180 50.940 -24.920 ;
        RECT 57.610 -25.200 57.870 -24.940 ;
        RECT 62.180 -25.160 62.440 -24.900 ;
        RECT 69.100 -25.200 69.360 -24.940 ;
        RECT 73.680 -25.200 73.940 -24.940 ;
        RECT 80.600 -25.230 80.860 -24.970 ;
        RECT 85.180 -25.210 85.440 -24.950 ;
        RECT 92.060 -25.210 92.360 -24.910 ;
        RECT -27.440 -25.660 -27.180 -25.400 ;
        RECT 135.320 -25.630 135.580 -25.370 ;
        RECT -15.650 -26.290 -15.390 -26.030 ;
        RECT 125.860 -26.130 126.120 -25.870 ;
        RECT 114.230 -26.630 114.490 -26.370 ;
        RECT -3.870 -27.040 -3.610 -26.780 ;
        RECT 102.100 -27.260 102.360 -27.000 ;
        RECT 8.110 -27.750 8.370 -27.490 ;
        RECT 90.360 -27.890 90.620 -27.630 ;
        RECT 19.780 -28.550 20.040 -28.290 ;
        RECT 78.480 -28.610 78.740 -28.350 ;
        RECT 31.370 -29.390 31.630 -29.130 ;
        RECT 66.460 -29.410 66.720 -29.150 ;
        RECT 43.110 -30.100 43.370 -29.840 ;
        RECT 54.960 -30.280 55.220 -30.020 ;
        RECT -39.880 -31.510 -39.620 -31.250 ;
        RECT -35.220 -33.870 -34.960 -33.610 ;
        RECT -23.720 -33.870 -23.460 -33.610 ;
        RECT -11.900 -33.870 -11.640 -33.610 ;
        RECT -0.090 -33.870 0.170 -33.610 ;
        RECT 11.720 -33.870 11.980 -33.610 ;
        RECT 23.540 -33.870 23.800 -33.610 ;
        RECT 35.360 -33.870 35.620 -33.610 ;
        RECT 47.180 -33.870 47.440 -33.610 ;
        RECT 59.000 -33.870 59.260 -33.610 ;
        RECT 70.820 -33.870 71.080 -33.610 ;
        RECT 82.640 -33.870 82.900 -33.610 ;
        RECT 94.480 -33.870 94.740 -33.610 ;
        RECT 106.320 -33.870 106.580 -33.610 ;
        RECT 118.190 -33.870 118.450 -33.610 ;
        RECT 130.060 -33.870 130.320 -33.610 ;
        RECT 139.070 -33.870 139.330 -33.610 ;
        RECT -31.480 -36.100 -31.220 -35.840 ;
        RECT -19.930 -36.100 -19.670 -35.840 ;
        RECT -8.240 -36.100 -7.980 -35.840 ;
        RECT 3.670 -36.100 3.930 -35.840 ;
        RECT 15.440 -36.100 15.700 -35.840 ;
        RECT 27.210 -36.100 27.470 -35.840 ;
        RECT 39.030 -36.100 39.290 -35.840 ;
        RECT 50.890 -36.100 51.150 -35.840 ;
        RECT 62.680 -36.100 62.940 -35.840 ;
        RECT 74.560 -36.100 74.820 -35.840 ;
        RECT 86.290 -36.100 86.550 -35.840 ;
        RECT 98.110 -36.100 98.370 -35.840 ;
        RECT 110.000 -36.100 110.260 -35.840 ;
        RECT 121.950 -36.100 122.210 -35.840 ;
        RECT 133.710 -36.100 133.970 -35.840 ;
        RECT 142.750 -36.100 143.010 -35.840 ;
        RECT -40.540 -36.540 -40.280 -36.280 ;
        RECT -41.200 -36.940 -40.940 -36.680 ;
        RECT -39.270 -41.630 -38.950 -41.310 ;
        RECT -27.430 -41.610 -27.170 -41.350 ;
        RECT -15.640 -41.610 -15.380 -41.350 ;
        RECT -3.860 -41.610 -3.600 -41.350 ;
        RECT 8.120 -41.610 8.380 -41.350 ;
        RECT 19.790 -41.600 20.050 -41.340 ;
        RECT 31.380 -41.590 31.640 -41.330 ;
        RECT 43.120 -41.590 43.380 -41.330 ;
        RECT 54.970 -41.590 55.230 -41.330 ;
        RECT 66.470 -41.610 66.730 -41.350 ;
        RECT 78.490 -41.610 78.750 -41.350 ;
        RECT 90.370 -41.610 90.630 -41.350 ;
        RECT 102.110 -41.610 102.370 -41.350 ;
        RECT 114.240 -41.600 114.500 -41.340 ;
        RECT 125.870 -41.610 126.130 -41.350 ;
        RECT 135.330 -41.600 135.590 -41.340 ;
        RECT -41.780 -43.720 -41.520 -43.460 ;
        RECT -39.130 -43.720 -38.870 -43.460 ;
        RECT -32.910 -43.720 -32.650 -43.460 ;
        RECT -21.410 -43.720 -21.150 -43.460 ;
        RECT -9.590 -43.720 -9.330 -43.460 ;
        RECT 2.220 -43.720 2.480 -43.460 ;
        RECT 14.030 -43.720 14.290 -43.460 ;
        RECT 25.850 -43.720 26.110 -43.460 ;
        RECT 37.670 -43.720 37.930 -43.460 ;
        RECT 49.490 -43.720 49.750 -43.460 ;
        RECT 61.310 -43.720 61.570 -43.460 ;
        RECT 73.130 -43.720 73.390 -43.460 ;
        RECT 84.950 -43.720 85.210 -43.460 ;
        RECT 96.790 -43.720 97.050 -43.460 ;
        RECT 108.630 -43.720 108.890 -43.460 ;
        RECT 120.500 -43.720 120.760 -43.460 ;
        RECT 132.370 -43.720 132.630 -43.460 ;
        RECT 141.380 -43.720 141.640 -43.460 ;
        RECT -37.870 -44.210 -37.610 -43.950 ;
        RECT -26.370 -44.210 -26.110 -43.950 ;
        RECT -14.550 -44.210 -14.290 -43.950 ;
        RECT -2.740 -44.210 -2.480 -43.950 ;
        RECT 9.070 -44.210 9.330 -43.950 ;
        RECT 20.890 -44.210 21.150 -43.950 ;
        RECT 32.710 -44.210 32.970 -43.950 ;
        RECT 44.530 -44.210 44.790 -43.950 ;
        RECT 56.350 -44.210 56.610 -43.950 ;
        RECT 68.170 -44.210 68.430 -43.950 ;
        RECT 79.990 -44.210 80.250 -43.950 ;
        RECT 91.830 -44.210 92.090 -43.950 ;
        RECT 103.670 -44.210 103.930 -43.950 ;
        RECT 115.540 -44.210 115.800 -43.950 ;
        RECT 127.410 -44.210 127.670 -43.950 ;
        RECT 136.420 -44.210 136.680 -43.950 ;
        RECT 144.460 -44.710 144.720 -44.450 ;
        RECT -32.870 -45.220 -32.610 -44.960 ;
        RECT -21.370 -45.220 -21.110 -44.960 ;
        RECT -9.550 -45.220 -9.290 -44.960 ;
        RECT 2.260 -45.220 2.520 -44.960 ;
        RECT 14.070 -45.220 14.330 -44.960 ;
        RECT 25.890 -45.220 26.150 -44.960 ;
        RECT 37.710 -45.220 37.970 -44.960 ;
        RECT 49.530 -45.220 49.790 -44.960 ;
        RECT 61.350 -45.220 61.610 -44.960 ;
        RECT 73.170 -45.220 73.430 -44.960 ;
        RECT 84.990 -45.220 85.250 -44.960 ;
        RECT 96.830 -45.220 97.090 -44.960 ;
        RECT 108.670 -45.220 108.930 -44.960 ;
        RECT 120.540 -45.220 120.800 -44.960 ;
        RECT 132.410 -45.220 132.670 -44.960 ;
        RECT 141.420 -45.220 141.680 -44.960 ;
        RECT 145.020 -45.600 145.280 -45.340 ;
        RECT -39.130 -46.620 -38.870 -46.360 ;
        RECT -32.910 -46.620 -32.650 -46.360 ;
        RECT -21.410 -46.620 -21.150 -46.360 ;
        RECT -9.590 -46.620 -9.330 -46.360 ;
        RECT 2.220 -46.620 2.480 -46.360 ;
        RECT 14.030 -46.620 14.290 -46.360 ;
        RECT 25.850 -46.620 26.110 -46.360 ;
        RECT 37.670 -46.620 37.930 -46.360 ;
        RECT 49.490 -46.620 49.750 -46.360 ;
        RECT 61.310 -46.620 61.570 -46.360 ;
        RECT 73.130 -46.620 73.390 -46.360 ;
        RECT 84.950 -46.620 85.210 -46.360 ;
        RECT 96.790 -46.620 97.050 -46.360 ;
        RECT 108.630 -46.620 108.890 -46.360 ;
        RECT 120.500 -46.620 120.760 -46.360 ;
        RECT 132.370 -46.620 132.630 -46.360 ;
        RECT 141.380 -46.620 141.640 -46.360 ;
        RECT -37.880 -48.750 -37.620 -48.490 ;
        RECT -26.380 -48.750 -26.120 -48.490 ;
        RECT -14.560 -48.750 -14.300 -48.490 ;
        RECT -2.750 -48.750 -2.490 -48.490 ;
        RECT 9.060 -48.750 9.320 -48.490 ;
        RECT 20.880 -48.750 21.140 -48.490 ;
        RECT 32.700 -48.750 32.960 -48.490 ;
        RECT 44.520 -48.750 44.780 -48.490 ;
        RECT 56.340 -48.750 56.600 -48.490 ;
        RECT 68.160 -48.750 68.420 -48.490 ;
        RECT 79.980 -48.750 80.240 -48.490 ;
        RECT 91.820 -48.750 92.080 -48.490 ;
        RECT 103.660 -48.750 103.920 -48.490 ;
        RECT 115.530 -48.750 115.790 -48.490 ;
        RECT 127.400 -48.750 127.660 -48.490 ;
        RECT 136.410 -48.750 136.670 -48.490 ;
        RECT -41.200 -53.400 -40.940 -53.140 ;
        RECT -40.540 -53.800 -40.280 -53.540 ;
        RECT -31.070 -54.230 -30.810 -53.970 ;
        RECT -19.530 -54.230 -19.270 -53.970 ;
        RECT -7.840 -54.230 -7.580 -53.970 ;
        RECT 4.070 -54.230 4.330 -53.970 ;
        RECT 15.840 -54.230 16.100 -53.970 ;
        RECT 27.610 -54.230 27.870 -53.970 ;
        RECT 39.430 -54.230 39.690 -53.970 ;
        RECT 51.290 -54.230 51.550 -53.970 ;
        RECT 63.080 -54.230 63.340 -53.970 ;
        RECT 74.960 -54.230 75.220 -53.970 ;
        RECT 86.690 -54.230 86.950 -53.970 ;
        RECT 98.510 -54.230 98.770 -53.970 ;
        RECT 110.400 -54.230 110.660 -53.970 ;
        RECT 122.350 -54.230 122.610 -53.970 ;
        RECT 134.110 -54.230 134.370 -53.970 ;
        RECT 143.150 -54.230 143.410 -53.970 ;
        RECT -35.220 -56.470 -34.960 -56.210 ;
        RECT -23.720 -56.470 -23.460 -56.210 ;
        RECT -11.900 -56.470 -11.640 -56.210 ;
        RECT -0.090 -56.470 0.170 -56.210 ;
        RECT 11.720 -56.470 11.980 -56.210 ;
        RECT 23.540 -56.470 23.800 -56.210 ;
        RECT 35.360 -56.470 35.620 -56.210 ;
        RECT 47.180 -56.470 47.440 -56.210 ;
        RECT 59.000 -56.470 59.260 -56.210 ;
        RECT 70.820 -56.470 71.080 -56.210 ;
        RECT 82.640 -56.470 82.900 -56.210 ;
        RECT 94.480 -56.470 94.740 -56.210 ;
        RECT 106.320 -56.470 106.580 -56.210 ;
        RECT 118.190 -56.470 118.450 -56.210 ;
        RECT 130.060 -56.470 130.320 -56.210 ;
        RECT 139.070 -56.470 139.330 -56.210 ;
        RECT -39.870 -58.830 -39.610 -58.570 ;
        RECT -35.220 -61.200 -34.960 -60.940 ;
        RECT -23.720 -61.200 -23.460 -60.940 ;
        RECT -11.900 -61.200 -11.640 -60.940 ;
        RECT -0.090 -61.200 0.170 -60.940 ;
        RECT 11.720 -61.200 11.980 -60.940 ;
        RECT 23.540 -61.200 23.800 -60.940 ;
        RECT 35.360 -61.200 35.620 -60.940 ;
        RECT 47.180 -61.200 47.440 -60.940 ;
        RECT 59.000 -61.200 59.260 -60.940 ;
        RECT 70.820 -61.200 71.080 -60.940 ;
        RECT 82.640 -61.200 82.900 -60.940 ;
        RECT 94.480 -61.200 94.740 -60.940 ;
        RECT 106.320 -61.200 106.580 -60.940 ;
        RECT 118.190 -61.200 118.450 -60.940 ;
        RECT 130.060 -61.200 130.320 -60.940 ;
        RECT 139.070 -61.200 139.330 -60.940 ;
        RECT -30.670 -63.430 -30.410 -63.170 ;
        RECT -19.110 -63.430 -18.850 -63.170 ;
        RECT -7.420 -63.430 -7.160 -63.170 ;
        RECT 4.490 -63.430 4.750 -63.170 ;
        RECT 16.260 -63.430 16.520 -63.170 ;
        RECT 28.030 -63.430 28.290 -63.170 ;
        RECT 39.850 -63.430 40.110 -63.170 ;
        RECT 51.710 -63.430 51.970 -63.170 ;
        RECT 63.500 -63.430 63.760 -63.170 ;
        RECT 75.380 -63.430 75.640 -63.170 ;
        RECT 87.110 -63.430 87.370 -63.170 ;
        RECT 98.930 -63.430 99.190 -63.170 ;
        RECT 110.820 -63.430 111.080 -63.170 ;
        RECT 122.770 -63.430 123.030 -63.170 ;
        RECT 134.530 -63.430 134.790 -63.170 ;
        RECT 143.570 -63.430 143.830 -63.170 ;
        RECT -40.540 -63.870 -40.280 -63.610 ;
        RECT -41.200 -64.270 -40.940 -64.010 ;
        RECT -37.870 -66.330 -37.610 -66.070 ;
        RECT -26.370 -66.330 -26.110 -66.070 ;
        RECT -14.550 -66.330 -14.290 -66.070 ;
        RECT -2.740 -66.330 -2.480 -66.070 ;
        RECT 9.070 -66.330 9.330 -66.070 ;
        RECT 20.890 -66.330 21.150 -66.070 ;
        RECT 32.710 -66.330 32.970 -66.070 ;
        RECT 44.530 -66.330 44.790 -66.070 ;
        RECT 56.350 -66.330 56.610 -66.070 ;
        RECT 68.170 -66.330 68.430 -66.070 ;
        RECT 79.990 -66.330 80.250 -66.070 ;
        RECT 91.830 -66.330 92.090 -66.070 ;
        RECT 103.670 -66.330 103.930 -66.070 ;
        RECT 115.540 -66.330 115.800 -66.070 ;
        RECT 127.410 -66.330 127.670 -66.070 ;
        RECT 136.420 -66.330 136.680 -66.070 ;
        RECT -37.880 -68.920 -37.620 -68.660 ;
        RECT -26.380 -68.920 -26.120 -68.660 ;
        RECT -14.560 -68.920 -14.300 -68.660 ;
        RECT -2.750 -68.920 -2.490 -68.660 ;
        RECT 9.060 -68.920 9.320 -68.660 ;
        RECT 20.880 -68.920 21.140 -68.660 ;
        RECT 32.700 -68.920 32.960 -68.660 ;
        RECT 44.520 -68.920 44.780 -68.660 ;
        RECT 56.340 -68.920 56.600 -68.660 ;
        RECT 68.160 -68.920 68.420 -68.660 ;
        RECT 79.980 -68.920 80.240 -68.660 ;
        RECT 91.820 -68.920 92.080 -68.660 ;
        RECT 103.660 -68.920 103.920 -68.660 ;
        RECT 115.530 -68.920 115.790 -68.660 ;
        RECT 127.400 -68.920 127.660 -68.660 ;
        RECT 136.410 -68.920 136.670 -68.660 ;
        RECT -39.130 -71.050 -38.870 -70.790 ;
        RECT -32.970 -71.050 -32.710 -70.790 ;
        RECT -21.470 -71.050 -21.210 -70.790 ;
        RECT -9.650 -71.050 -9.390 -70.790 ;
        RECT 2.160 -71.050 2.420 -70.790 ;
        RECT 13.970 -71.050 14.230 -70.790 ;
        RECT 25.790 -71.050 26.050 -70.790 ;
        RECT 37.610 -71.050 37.870 -70.790 ;
        RECT 49.430 -71.050 49.690 -70.790 ;
        RECT 61.250 -71.050 61.510 -70.790 ;
        RECT 73.070 -71.050 73.330 -70.790 ;
        RECT 84.890 -71.050 85.150 -70.790 ;
        RECT 96.730 -71.050 96.990 -70.790 ;
        RECT 108.570 -71.050 108.830 -70.790 ;
        RECT 120.440 -71.050 120.700 -70.790 ;
        RECT 132.310 -71.050 132.570 -70.790 ;
        RECT 141.320 -71.050 141.580 -70.790 ;
        RECT 145.560 -71.970 145.820 -71.710 ;
        RECT -32.910 -72.560 -32.650 -72.300 ;
        RECT -21.410 -72.560 -21.150 -72.300 ;
        RECT -9.590 -72.560 -9.330 -72.300 ;
        RECT 2.220 -72.560 2.480 -72.300 ;
        RECT 14.030 -72.560 14.290 -72.300 ;
        RECT 25.850 -72.560 26.110 -72.300 ;
        RECT 37.670 -72.560 37.930 -72.300 ;
        RECT 49.490 -72.560 49.750 -72.300 ;
        RECT 61.310 -72.560 61.570 -72.300 ;
        RECT 73.130 -72.560 73.390 -72.300 ;
        RECT 84.950 -72.560 85.210 -72.300 ;
        RECT 96.790 -72.560 97.050 -72.300 ;
        RECT 108.630 -72.560 108.890 -72.300 ;
        RECT 120.500 -72.560 120.760 -72.300 ;
        RECT 132.370 -72.560 132.630 -72.300 ;
        RECT 141.380 -72.560 141.640 -72.300 ;
        RECT 146.110 -72.940 146.370 -72.680 ;
        RECT -39.130 -73.950 -38.870 -73.690 ;
        RECT -32.970 -73.950 -32.710 -73.690 ;
        RECT -21.470 -73.950 -21.210 -73.690 ;
        RECT -9.650 -73.950 -9.390 -73.690 ;
        RECT 2.160 -73.950 2.420 -73.690 ;
        RECT 13.970 -73.950 14.230 -73.690 ;
        RECT 25.790 -73.950 26.050 -73.690 ;
        RECT 37.610 -73.950 37.870 -73.690 ;
        RECT 49.430 -73.950 49.690 -73.690 ;
        RECT 61.250 -73.950 61.510 -73.690 ;
        RECT 73.070 -73.950 73.330 -73.690 ;
        RECT 84.890 -73.950 85.150 -73.690 ;
        RECT 96.730 -73.950 96.990 -73.690 ;
        RECT 108.570 -73.950 108.830 -73.690 ;
        RECT 120.440 -73.950 120.700 -73.690 ;
        RECT 132.310 -73.950 132.570 -73.690 ;
        RECT 141.320 -73.950 141.580 -73.690 ;
        RECT -37.880 -76.090 -37.620 -75.830 ;
        RECT -26.380 -76.090 -26.120 -75.830 ;
        RECT -14.560 -76.090 -14.300 -75.830 ;
        RECT -2.750 -76.090 -2.490 -75.830 ;
        RECT 9.060 -76.090 9.320 -75.830 ;
        RECT 20.880 -76.090 21.140 -75.830 ;
        RECT 32.700 -76.090 32.960 -75.830 ;
        RECT 44.520 -76.090 44.780 -75.830 ;
        RECT 56.340 -76.090 56.600 -75.830 ;
        RECT 68.160 -76.090 68.420 -75.830 ;
        RECT 79.980 -76.090 80.240 -75.830 ;
        RECT 91.820 -76.090 92.080 -75.830 ;
        RECT 103.660 -76.090 103.920 -75.830 ;
        RECT 115.530 -76.090 115.790 -75.830 ;
        RECT 127.400 -76.090 127.660 -75.830 ;
        RECT 136.410 -76.090 136.670 -75.830 ;
        RECT -41.200 -80.730 -40.940 -80.470 ;
        RECT -40.540 -81.130 -40.280 -80.870 ;
        RECT -30.260 -81.560 -30.000 -81.300 ;
        RECT -18.700 -81.560 -18.440 -81.300 ;
        RECT -7.010 -81.560 -6.750 -81.300 ;
        RECT 4.900 -81.560 5.160 -81.300 ;
        RECT 16.670 -81.560 16.930 -81.300 ;
        RECT 28.440 -81.560 28.700 -81.300 ;
        RECT 40.260 -81.560 40.520 -81.300 ;
        RECT 52.120 -81.560 52.380 -81.300 ;
        RECT 63.910 -81.560 64.170 -81.300 ;
        RECT 75.790 -81.560 76.050 -81.300 ;
        RECT 87.520 -81.560 87.780 -81.300 ;
        RECT 99.340 -81.560 99.600 -81.300 ;
        RECT 111.230 -81.560 111.490 -81.300 ;
        RECT 123.180 -81.560 123.440 -81.300 ;
        RECT 134.940 -81.560 135.200 -81.300 ;
        RECT 143.980 -81.560 144.240 -81.300 ;
        RECT -35.220 -83.800 -34.960 -83.540 ;
        RECT -23.720 -83.800 -23.460 -83.540 ;
        RECT -11.900 -83.800 -11.640 -83.540 ;
        RECT -0.090 -83.800 0.170 -83.540 ;
        RECT 11.720 -83.800 11.980 -83.540 ;
        RECT 23.540 -83.800 23.800 -83.540 ;
        RECT 35.360 -83.800 35.620 -83.540 ;
        RECT 47.180 -83.800 47.440 -83.540 ;
        RECT 59.000 -83.800 59.260 -83.540 ;
        RECT 70.820 -83.800 71.080 -83.540 ;
        RECT 82.640 -83.800 82.900 -83.540 ;
        RECT 94.480 -83.800 94.740 -83.540 ;
        RECT 106.320 -83.800 106.580 -83.540 ;
        RECT 118.190 -83.800 118.450 -83.540 ;
        RECT 130.060 -83.800 130.320 -83.540 ;
        RECT 139.070 -83.800 139.330 -83.540 ;
        RECT -39.880 -86.160 -39.620 -85.900 ;
      LAYER met2 ;
        RECT -43.140 50.260 -42.840 50.660 ;
        RECT -43.060 -30.580 -42.920 50.260 ;
        RECT 1.290 48.350 1.550 48.670 ;
        RECT 1.350 47.840 1.500 48.350 ;
        RECT 3.050 48.290 3.190 50.590 ;
        RECT 3.960 49.750 4.100 50.590 ;
        RECT 5.190 50.340 5.590 50.740 ;
        RECT 3.960 49.330 4.350 49.750 ;
        RECT 5.320 49.720 5.460 50.340 ;
        RECT 6.660 49.750 6.800 50.590 ;
        RECT 5.230 49.400 5.550 49.720 ;
        RECT 3.960 48.290 4.100 49.330 ;
        RECT 2.960 47.980 3.280 48.290 ;
        RECT 3.870 47.980 4.190 48.290 ;
        RECT 5.320 48.200 5.460 49.400 ;
        RECT 6.400 49.330 6.800 49.750 ;
        RECT 1.250 47.520 1.570 47.840 ;
        RECT 1.350 46.980 1.500 47.520 ;
        RECT 1.270 46.660 1.590 46.980 ;
        RECT 1.350 46.260 1.500 46.660 ;
        RECT 1.280 45.940 1.540 46.260 ;
        RECT 1.350 45.410 1.500 45.940 ;
        RECT 3.050 45.880 3.190 47.980 ;
        RECT 3.960 45.880 4.100 47.980 ;
        RECT 5.320 47.890 5.830 48.200 ;
        RECT 5.320 46.620 5.460 47.890 ;
        RECT 6.660 46.620 6.800 49.330 ;
        RECT 7.580 46.620 7.720 50.590 ;
        RECT 8.800 48.290 8.940 50.590 ;
        RECT 9.710 49.750 9.850 50.590 ;
        RECT 10.950 50.340 11.350 50.740 ;
        RECT 9.710 49.330 10.100 49.750 ;
        RECT 11.070 49.720 11.210 50.340 ;
        RECT 12.410 49.750 12.550 50.590 ;
        RECT 10.980 49.400 11.300 49.720 ;
        RECT 9.710 48.290 9.850 49.330 ;
        RECT 8.710 47.980 9.030 48.290 ;
        RECT 9.620 47.980 9.940 48.290 ;
        RECT 11.070 48.200 11.210 49.400 ;
        RECT 12.150 49.330 12.550 49.750 ;
        RECT 4.930 46.310 5.460 46.620 ;
        RECT 6.570 46.310 6.890 46.620 ;
        RECT 7.480 46.310 7.800 46.620 ;
        RECT 2.960 45.570 3.280 45.880 ;
        RECT 3.870 45.570 4.190 45.880 ;
        RECT 5.320 45.790 5.460 46.310 ;
        RECT 1.260 45.090 1.580 45.410 ;
        RECT 1.350 44.610 1.500 45.090 ;
        RECT 1.260 44.290 1.580 44.610 ;
        RECT 1.350 43.850 1.500 44.290 ;
        RECT 1.280 43.530 1.540 43.850 ;
        RECT 1.350 42.480 1.500 43.530 ;
        RECT 3.050 42.910 3.190 45.570 ;
        RECT 3.960 42.910 4.100 45.570 ;
        RECT 5.320 45.480 5.830 45.790 ;
        RECT 5.320 44.210 5.460 45.480 ;
        RECT 6.660 44.210 6.800 46.310 ;
        RECT 7.580 44.210 7.720 46.310 ;
        RECT 8.800 45.880 8.940 47.980 ;
        RECT 9.710 45.880 9.850 47.980 ;
        RECT 11.070 47.890 11.580 48.200 ;
        RECT 11.070 46.620 11.210 47.890 ;
        RECT 12.410 46.620 12.550 49.330 ;
        RECT 13.330 46.620 13.470 50.590 ;
        RECT 14.550 48.290 14.690 50.590 ;
        RECT 15.460 49.750 15.600 50.590 ;
        RECT 16.700 50.340 17.100 50.740 ;
        RECT 15.460 49.330 15.850 49.750 ;
        RECT 16.820 49.720 16.960 50.340 ;
        RECT 18.160 49.750 18.300 50.590 ;
        RECT 16.730 49.400 17.050 49.720 ;
        RECT 15.460 48.290 15.600 49.330 ;
        RECT 14.460 47.980 14.780 48.290 ;
        RECT 15.370 47.980 15.690 48.290 ;
        RECT 16.820 48.200 16.960 49.400 ;
        RECT 17.900 49.330 18.300 49.750 ;
        RECT 10.680 46.310 11.210 46.620 ;
        RECT 12.320 46.310 12.640 46.620 ;
        RECT 13.230 46.310 13.550 46.620 ;
        RECT 8.710 45.570 9.030 45.880 ;
        RECT 9.620 45.570 9.940 45.880 ;
        RECT 11.070 45.790 11.210 46.310 ;
        RECT 4.930 43.900 5.460 44.210 ;
        RECT 6.570 43.900 6.890 44.210 ;
        RECT 7.480 43.900 7.800 44.210 ;
        RECT 2.960 42.600 3.280 42.910 ;
        RECT 3.870 42.600 4.190 42.910 ;
        RECT 5.320 42.820 5.460 43.900 ;
        RECT 1.270 42.160 1.590 42.480 ;
        RECT 1.350 41.620 1.500 42.160 ;
        RECT 1.270 41.300 1.590 41.620 ;
        RECT 1.350 40.880 1.500 41.300 ;
        RECT 1.280 40.560 1.540 40.880 ;
        RECT 1.350 40.050 1.500 40.560 ;
        RECT 3.050 40.500 3.190 42.600 ;
        RECT 3.960 40.500 4.100 42.600 ;
        RECT 5.320 42.510 5.830 42.820 ;
        RECT 5.320 41.240 5.460 42.510 ;
        RECT 6.660 41.240 6.800 43.900 ;
        RECT 7.580 41.240 7.720 43.900 ;
        RECT 8.800 42.910 8.940 45.570 ;
        RECT 9.710 42.910 9.850 45.570 ;
        RECT 11.070 45.480 11.580 45.790 ;
        RECT 11.070 44.210 11.210 45.480 ;
        RECT 12.410 44.210 12.550 46.310 ;
        RECT 13.330 44.210 13.470 46.310 ;
        RECT 14.550 45.880 14.690 47.980 ;
        RECT 15.460 45.880 15.600 47.980 ;
        RECT 16.820 47.890 17.330 48.200 ;
        RECT 16.820 46.620 16.960 47.890 ;
        RECT 18.160 46.620 18.300 49.330 ;
        RECT 19.080 46.620 19.220 50.590 ;
        RECT 20.300 48.290 20.440 50.590 ;
        RECT 21.210 49.750 21.350 50.590 ;
        RECT 22.430 50.340 22.830 50.740 ;
        RECT 21.210 49.330 21.600 49.750 ;
        RECT 22.570 49.720 22.710 50.340 ;
        RECT 23.910 49.750 24.050 50.590 ;
        RECT 22.480 49.400 22.800 49.720 ;
        RECT 21.210 48.290 21.350 49.330 ;
        RECT 20.210 47.980 20.530 48.290 ;
        RECT 21.120 47.980 21.440 48.290 ;
        RECT 22.570 48.200 22.710 49.400 ;
        RECT 23.650 49.330 24.050 49.750 ;
        RECT 16.430 46.310 16.960 46.620 ;
        RECT 18.070 46.310 18.390 46.620 ;
        RECT 18.980 46.310 19.300 46.620 ;
        RECT 14.460 45.570 14.780 45.880 ;
        RECT 15.370 45.570 15.690 45.880 ;
        RECT 16.820 45.790 16.960 46.310 ;
        RECT 10.680 43.900 11.210 44.210 ;
        RECT 12.320 43.900 12.640 44.210 ;
        RECT 13.230 43.900 13.550 44.210 ;
        RECT 8.710 42.600 9.030 42.910 ;
        RECT 9.620 42.600 9.940 42.910 ;
        RECT 11.070 42.820 11.210 43.900 ;
        RECT 4.930 40.930 5.460 41.240 ;
        RECT 6.570 40.930 6.890 41.240 ;
        RECT 7.480 40.930 7.800 41.240 ;
        RECT 2.960 40.190 3.280 40.500 ;
        RECT 3.870 40.190 4.190 40.500 ;
        RECT 5.320 40.410 5.460 40.930 ;
        RECT 1.270 39.730 1.590 40.050 ;
        RECT 1.350 39.210 1.500 39.730 ;
        RECT 1.270 38.890 1.590 39.210 ;
        RECT 1.350 38.470 1.500 38.890 ;
        RECT 1.290 38.150 1.550 38.470 ;
        RECT 1.350 36.060 1.500 38.150 ;
        RECT 3.050 38.090 3.190 40.190 ;
        RECT 3.960 38.090 4.100 40.190 ;
        RECT 5.320 40.100 5.830 40.410 ;
        RECT 5.320 38.830 5.460 40.100 ;
        RECT 6.660 38.830 6.800 40.930 ;
        RECT 7.580 38.830 7.720 40.930 ;
        RECT 8.800 40.500 8.940 42.600 ;
        RECT 9.710 40.500 9.850 42.600 ;
        RECT 11.070 42.510 11.580 42.820 ;
        RECT 11.070 41.240 11.210 42.510 ;
        RECT 12.410 41.240 12.550 43.900 ;
        RECT 13.330 41.240 13.470 43.900 ;
        RECT 14.550 42.910 14.690 45.570 ;
        RECT 15.460 42.910 15.600 45.570 ;
        RECT 16.820 45.480 17.330 45.790 ;
        RECT 16.820 44.210 16.960 45.480 ;
        RECT 18.160 44.210 18.300 46.310 ;
        RECT 19.080 44.210 19.220 46.310 ;
        RECT 20.300 45.880 20.440 47.980 ;
        RECT 21.210 45.880 21.350 47.980 ;
        RECT 22.570 47.890 23.080 48.200 ;
        RECT 22.570 46.620 22.710 47.890 ;
        RECT 23.910 46.620 24.050 49.330 ;
        RECT 24.830 46.620 24.970 50.590 ;
        RECT 26.050 48.290 26.190 50.590 ;
        RECT 26.960 49.750 27.100 50.590 ;
        RECT 28.190 50.340 28.590 50.740 ;
        RECT 26.960 49.330 27.350 49.750 ;
        RECT 28.320 49.720 28.460 50.340 ;
        RECT 29.660 49.750 29.800 50.590 ;
        RECT 28.230 49.400 28.550 49.720 ;
        RECT 26.960 48.290 27.100 49.330 ;
        RECT 25.960 47.980 26.280 48.290 ;
        RECT 26.870 47.980 27.190 48.290 ;
        RECT 28.320 48.200 28.460 49.400 ;
        RECT 29.400 49.330 29.800 49.750 ;
        RECT 22.180 46.310 22.710 46.620 ;
        RECT 23.820 46.310 24.140 46.620 ;
        RECT 24.730 46.310 25.050 46.620 ;
        RECT 20.210 45.570 20.530 45.880 ;
        RECT 21.120 45.570 21.440 45.880 ;
        RECT 22.570 45.790 22.710 46.310 ;
        RECT 16.430 43.900 16.960 44.210 ;
        RECT 18.070 43.900 18.390 44.210 ;
        RECT 18.980 43.900 19.300 44.210 ;
        RECT 14.460 42.600 14.780 42.910 ;
        RECT 15.370 42.600 15.690 42.910 ;
        RECT 16.820 42.820 16.960 43.900 ;
        RECT 10.680 40.930 11.210 41.240 ;
        RECT 12.320 40.930 12.640 41.240 ;
        RECT 13.230 40.930 13.550 41.240 ;
        RECT 8.710 40.190 9.030 40.500 ;
        RECT 9.620 40.190 9.940 40.500 ;
        RECT 11.070 40.410 11.210 40.930 ;
        RECT 4.930 38.520 5.460 38.830 ;
        RECT 6.570 38.520 6.890 38.830 ;
        RECT 7.480 38.520 7.800 38.830 ;
        RECT 2.960 37.780 3.280 38.090 ;
        RECT 3.870 37.780 4.190 38.090 ;
        RECT 5.320 38.000 5.460 38.520 ;
        RECT 1.290 35.740 1.550 36.060 ;
        RECT 1.350 33.650 1.500 35.740 ;
        RECT 3.050 35.680 3.190 37.780 ;
        RECT 3.960 35.680 4.100 37.780 ;
        RECT 5.320 37.690 5.830 38.000 ;
        RECT 5.320 36.420 5.460 37.690 ;
        RECT 6.660 36.420 6.800 38.520 ;
        RECT 7.580 36.420 7.720 38.520 ;
        RECT 8.800 38.090 8.940 40.190 ;
        RECT 9.710 38.090 9.850 40.190 ;
        RECT 11.070 40.100 11.580 40.410 ;
        RECT 11.070 38.830 11.210 40.100 ;
        RECT 12.410 38.830 12.550 40.930 ;
        RECT 13.330 38.830 13.470 40.930 ;
        RECT 14.550 40.500 14.690 42.600 ;
        RECT 15.460 40.500 15.600 42.600 ;
        RECT 16.820 42.510 17.330 42.820 ;
        RECT 16.820 41.240 16.960 42.510 ;
        RECT 18.160 41.240 18.300 43.900 ;
        RECT 19.080 41.240 19.220 43.900 ;
        RECT 20.300 42.910 20.440 45.570 ;
        RECT 21.210 42.910 21.350 45.570 ;
        RECT 22.570 45.480 23.080 45.790 ;
        RECT 22.570 44.210 22.710 45.480 ;
        RECT 23.910 44.210 24.050 46.310 ;
        RECT 24.830 44.210 24.970 46.310 ;
        RECT 26.050 45.880 26.190 47.980 ;
        RECT 26.960 45.880 27.100 47.980 ;
        RECT 28.320 47.890 28.830 48.200 ;
        RECT 28.320 46.620 28.460 47.890 ;
        RECT 29.660 46.620 29.800 49.330 ;
        RECT 30.580 46.620 30.720 50.590 ;
        RECT 31.800 48.290 31.940 50.590 ;
        RECT 32.710 49.750 32.850 50.590 ;
        RECT 33.930 50.340 34.330 50.740 ;
        RECT 32.710 49.330 33.100 49.750 ;
        RECT 34.070 49.720 34.210 50.340 ;
        RECT 35.410 49.750 35.550 50.590 ;
        RECT 33.980 49.400 34.300 49.720 ;
        RECT 32.710 48.290 32.850 49.330 ;
        RECT 31.710 47.980 32.030 48.290 ;
        RECT 32.620 47.980 32.940 48.290 ;
        RECT 34.070 48.200 34.210 49.400 ;
        RECT 35.150 49.330 35.550 49.750 ;
        RECT 27.930 46.310 28.460 46.620 ;
        RECT 29.570 46.310 29.890 46.620 ;
        RECT 30.480 46.310 30.800 46.620 ;
        RECT 25.960 45.570 26.280 45.880 ;
        RECT 26.870 45.570 27.190 45.880 ;
        RECT 28.320 45.790 28.460 46.310 ;
        RECT 22.180 43.900 22.710 44.210 ;
        RECT 23.820 43.900 24.140 44.210 ;
        RECT 24.730 43.900 25.050 44.210 ;
        RECT 20.210 42.600 20.530 42.910 ;
        RECT 21.120 42.600 21.440 42.910 ;
        RECT 22.570 42.820 22.710 43.900 ;
        RECT 16.430 40.930 16.960 41.240 ;
        RECT 18.070 40.930 18.390 41.240 ;
        RECT 18.980 40.930 19.300 41.240 ;
        RECT 14.460 40.190 14.780 40.500 ;
        RECT 15.370 40.190 15.690 40.500 ;
        RECT 16.820 40.410 16.960 40.930 ;
        RECT 10.680 38.520 11.210 38.830 ;
        RECT 12.320 38.520 12.640 38.830 ;
        RECT 13.230 38.520 13.550 38.830 ;
        RECT 8.710 37.780 9.030 38.090 ;
        RECT 9.620 37.780 9.940 38.090 ;
        RECT 11.070 38.000 11.210 38.520 ;
        RECT 4.930 36.110 5.460 36.420 ;
        RECT 6.570 36.110 6.890 36.420 ;
        RECT 7.480 36.110 7.800 36.420 ;
        RECT 2.960 35.370 3.280 35.680 ;
        RECT 3.870 35.370 4.190 35.680 ;
        RECT 5.320 35.590 5.460 36.110 ;
        RECT 1.290 33.330 1.550 33.650 ;
        RECT 1.350 31.240 1.500 33.330 ;
        RECT 3.050 33.270 3.190 35.370 ;
        RECT 3.960 33.270 4.100 35.370 ;
        RECT 5.320 35.280 5.830 35.590 ;
        RECT 5.320 34.010 5.460 35.280 ;
        RECT 6.660 34.010 6.800 36.110 ;
        RECT 7.580 34.010 7.720 36.110 ;
        RECT 8.800 35.680 8.940 37.780 ;
        RECT 9.710 35.680 9.850 37.780 ;
        RECT 11.070 37.690 11.580 38.000 ;
        RECT 11.070 36.420 11.210 37.690 ;
        RECT 12.410 36.420 12.550 38.520 ;
        RECT 13.330 36.420 13.470 38.520 ;
        RECT 14.550 38.090 14.690 40.190 ;
        RECT 15.460 38.090 15.600 40.190 ;
        RECT 16.820 40.100 17.330 40.410 ;
        RECT 16.820 38.830 16.960 40.100 ;
        RECT 18.160 38.830 18.300 40.930 ;
        RECT 19.080 38.830 19.220 40.930 ;
        RECT 20.300 40.500 20.440 42.600 ;
        RECT 21.210 40.500 21.350 42.600 ;
        RECT 22.570 42.510 23.080 42.820 ;
        RECT 22.570 41.240 22.710 42.510 ;
        RECT 23.910 41.240 24.050 43.900 ;
        RECT 24.830 41.240 24.970 43.900 ;
        RECT 26.050 42.910 26.190 45.570 ;
        RECT 26.960 42.910 27.100 45.570 ;
        RECT 28.320 45.480 28.830 45.790 ;
        RECT 28.320 44.210 28.460 45.480 ;
        RECT 29.660 44.210 29.800 46.310 ;
        RECT 30.580 44.210 30.720 46.310 ;
        RECT 31.800 45.880 31.940 47.980 ;
        RECT 32.710 45.880 32.850 47.980 ;
        RECT 34.070 47.890 34.580 48.200 ;
        RECT 34.070 46.620 34.210 47.890 ;
        RECT 35.410 46.620 35.550 49.330 ;
        RECT 36.330 46.620 36.470 50.590 ;
        RECT 37.550 48.290 37.690 50.590 ;
        RECT 38.460 49.750 38.600 50.590 ;
        RECT 39.680 50.340 40.080 50.740 ;
        RECT 38.460 49.330 38.850 49.750 ;
        RECT 39.820 49.720 39.960 50.340 ;
        RECT 41.160 49.750 41.300 50.590 ;
        RECT 39.730 49.400 40.050 49.720 ;
        RECT 38.460 48.290 38.600 49.330 ;
        RECT 37.460 47.980 37.780 48.290 ;
        RECT 38.370 47.980 38.690 48.290 ;
        RECT 39.820 48.200 39.960 49.400 ;
        RECT 40.900 49.330 41.300 49.750 ;
        RECT 33.680 46.310 34.210 46.620 ;
        RECT 35.320 46.310 35.640 46.620 ;
        RECT 36.230 46.310 36.550 46.620 ;
        RECT 31.710 45.570 32.030 45.880 ;
        RECT 32.620 45.570 32.940 45.880 ;
        RECT 34.070 45.790 34.210 46.310 ;
        RECT 27.930 43.900 28.460 44.210 ;
        RECT 29.570 43.900 29.890 44.210 ;
        RECT 30.480 43.900 30.800 44.210 ;
        RECT 25.960 42.600 26.280 42.910 ;
        RECT 26.870 42.600 27.190 42.910 ;
        RECT 28.320 42.820 28.460 43.900 ;
        RECT 22.180 40.930 22.710 41.240 ;
        RECT 23.820 40.930 24.140 41.240 ;
        RECT 24.730 40.930 25.050 41.240 ;
        RECT 20.210 40.190 20.530 40.500 ;
        RECT 21.120 40.190 21.440 40.500 ;
        RECT 22.570 40.410 22.710 40.930 ;
        RECT 16.430 38.520 16.960 38.830 ;
        RECT 18.070 38.520 18.390 38.830 ;
        RECT 18.980 38.520 19.300 38.830 ;
        RECT 14.460 37.780 14.780 38.090 ;
        RECT 15.370 37.780 15.690 38.090 ;
        RECT 16.820 38.000 16.960 38.520 ;
        RECT 10.680 36.110 11.210 36.420 ;
        RECT 12.320 36.110 12.640 36.420 ;
        RECT 13.230 36.110 13.550 36.420 ;
        RECT 8.710 35.370 9.030 35.680 ;
        RECT 9.620 35.370 9.940 35.680 ;
        RECT 11.070 35.590 11.210 36.110 ;
        RECT 4.930 33.700 5.460 34.010 ;
        RECT 6.570 33.700 6.890 34.010 ;
        RECT 7.480 33.700 7.800 34.010 ;
        RECT 2.960 32.960 3.280 33.270 ;
        RECT 3.870 32.960 4.190 33.270 ;
        RECT 5.320 33.180 5.460 33.700 ;
        RECT 1.290 30.920 1.550 31.240 ;
        RECT 1.350 28.830 1.500 30.920 ;
        RECT 3.050 30.860 3.190 32.960 ;
        RECT 3.960 30.860 4.100 32.960 ;
        RECT 5.320 32.870 5.830 33.180 ;
        RECT 5.320 31.600 5.460 32.870 ;
        RECT 6.660 31.600 6.800 33.700 ;
        RECT 7.580 31.600 7.720 33.700 ;
        RECT 8.800 33.270 8.940 35.370 ;
        RECT 9.710 33.270 9.850 35.370 ;
        RECT 11.070 35.280 11.580 35.590 ;
        RECT 11.070 34.010 11.210 35.280 ;
        RECT 12.410 34.010 12.550 36.110 ;
        RECT 13.330 34.010 13.470 36.110 ;
        RECT 14.550 35.680 14.690 37.780 ;
        RECT 15.460 35.680 15.600 37.780 ;
        RECT 16.820 37.690 17.330 38.000 ;
        RECT 16.820 36.420 16.960 37.690 ;
        RECT 18.160 36.420 18.300 38.520 ;
        RECT 19.080 36.420 19.220 38.520 ;
        RECT 20.300 38.090 20.440 40.190 ;
        RECT 21.210 38.090 21.350 40.190 ;
        RECT 22.570 40.100 23.080 40.410 ;
        RECT 22.570 38.830 22.710 40.100 ;
        RECT 23.910 38.830 24.050 40.930 ;
        RECT 24.830 38.830 24.970 40.930 ;
        RECT 26.050 40.500 26.190 42.600 ;
        RECT 26.960 40.500 27.100 42.600 ;
        RECT 28.320 42.510 28.830 42.820 ;
        RECT 28.320 41.240 28.460 42.510 ;
        RECT 29.660 41.240 29.800 43.900 ;
        RECT 30.580 41.240 30.720 43.900 ;
        RECT 31.800 42.910 31.940 45.570 ;
        RECT 32.710 42.910 32.850 45.570 ;
        RECT 34.070 45.480 34.580 45.790 ;
        RECT 34.070 44.210 34.210 45.480 ;
        RECT 35.410 44.210 35.550 46.310 ;
        RECT 36.330 44.210 36.470 46.310 ;
        RECT 37.550 45.880 37.690 47.980 ;
        RECT 38.460 45.880 38.600 47.980 ;
        RECT 39.820 47.890 40.330 48.200 ;
        RECT 39.820 46.620 39.960 47.890 ;
        RECT 41.160 46.620 41.300 49.330 ;
        RECT 42.080 46.620 42.220 50.590 ;
        RECT 43.300 48.290 43.440 50.590 ;
        RECT 44.210 49.750 44.350 50.590 ;
        RECT 45.430 50.340 45.830 50.740 ;
        RECT 44.210 49.330 44.600 49.750 ;
        RECT 45.570 49.720 45.710 50.340 ;
        RECT 46.910 49.750 47.050 50.590 ;
        RECT 45.480 49.400 45.800 49.720 ;
        RECT 44.210 48.290 44.350 49.330 ;
        RECT 43.210 47.980 43.530 48.290 ;
        RECT 44.120 47.980 44.440 48.290 ;
        RECT 45.570 48.200 45.710 49.400 ;
        RECT 46.650 49.330 47.050 49.750 ;
        RECT 39.430 46.310 39.960 46.620 ;
        RECT 41.070 46.310 41.390 46.620 ;
        RECT 41.980 46.310 42.300 46.620 ;
        RECT 37.460 45.570 37.780 45.880 ;
        RECT 38.370 45.570 38.690 45.880 ;
        RECT 39.820 45.790 39.960 46.310 ;
        RECT 33.680 43.900 34.210 44.210 ;
        RECT 35.320 43.900 35.640 44.210 ;
        RECT 36.230 43.900 36.550 44.210 ;
        RECT 31.710 42.600 32.030 42.910 ;
        RECT 32.620 42.600 32.940 42.910 ;
        RECT 34.070 42.820 34.210 43.900 ;
        RECT 27.930 40.930 28.460 41.240 ;
        RECT 29.570 40.930 29.890 41.240 ;
        RECT 30.480 40.930 30.800 41.240 ;
        RECT 25.960 40.190 26.280 40.500 ;
        RECT 26.870 40.190 27.190 40.500 ;
        RECT 28.320 40.410 28.460 40.930 ;
        RECT 22.180 38.520 22.710 38.830 ;
        RECT 23.820 38.520 24.140 38.830 ;
        RECT 24.730 38.520 25.050 38.830 ;
        RECT 20.210 37.780 20.530 38.090 ;
        RECT 21.120 37.780 21.440 38.090 ;
        RECT 22.570 38.000 22.710 38.520 ;
        RECT 16.430 36.110 16.960 36.420 ;
        RECT 18.070 36.110 18.390 36.420 ;
        RECT 18.980 36.110 19.300 36.420 ;
        RECT 14.460 35.370 14.780 35.680 ;
        RECT 15.370 35.370 15.690 35.680 ;
        RECT 16.820 35.590 16.960 36.110 ;
        RECT 10.680 33.700 11.210 34.010 ;
        RECT 12.320 33.700 12.640 34.010 ;
        RECT 13.230 33.700 13.550 34.010 ;
        RECT 8.710 32.960 9.030 33.270 ;
        RECT 9.620 32.960 9.940 33.270 ;
        RECT 11.070 33.180 11.210 33.700 ;
        RECT 4.930 31.290 5.460 31.600 ;
        RECT 6.570 31.290 6.890 31.600 ;
        RECT 7.480 31.290 7.800 31.600 ;
        RECT 2.960 30.550 3.280 30.860 ;
        RECT 3.870 30.550 4.190 30.860 ;
        RECT 5.320 30.770 5.460 31.290 ;
        RECT 1.290 28.510 1.550 28.830 ;
        RECT 1.350 26.020 1.500 28.510 ;
        RECT 3.050 28.050 3.190 30.550 ;
        RECT 3.960 28.050 4.100 30.550 ;
        RECT 5.320 30.460 5.830 30.770 ;
        RECT 5.320 29.190 5.460 30.460 ;
        RECT 6.660 29.190 6.800 31.290 ;
        RECT 7.580 29.190 7.720 31.290 ;
        RECT 8.800 30.860 8.940 32.960 ;
        RECT 9.710 30.860 9.850 32.960 ;
        RECT 11.070 32.870 11.580 33.180 ;
        RECT 11.070 31.600 11.210 32.870 ;
        RECT 12.410 31.600 12.550 33.700 ;
        RECT 13.330 31.600 13.470 33.700 ;
        RECT 14.550 33.270 14.690 35.370 ;
        RECT 15.460 33.270 15.600 35.370 ;
        RECT 16.820 35.280 17.330 35.590 ;
        RECT 16.820 34.010 16.960 35.280 ;
        RECT 18.160 34.010 18.300 36.110 ;
        RECT 19.080 34.010 19.220 36.110 ;
        RECT 20.300 35.680 20.440 37.780 ;
        RECT 21.210 35.680 21.350 37.780 ;
        RECT 22.570 37.690 23.080 38.000 ;
        RECT 22.570 36.420 22.710 37.690 ;
        RECT 23.910 36.420 24.050 38.520 ;
        RECT 24.830 36.420 24.970 38.520 ;
        RECT 26.050 38.090 26.190 40.190 ;
        RECT 26.960 38.090 27.100 40.190 ;
        RECT 28.320 40.100 28.830 40.410 ;
        RECT 28.320 38.830 28.460 40.100 ;
        RECT 29.660 38.830 29.800 40.930 ;
        RECT 30.580 38.830 30.720 40.930 ;
        RECT 31.800 40.500 31.940 42.600 ;
        RECT 32.710 40.500 32.850 42.600 ;
        RECT 34.070 42.510 34.580 42.820 ;
        RECT 34.070 41.240 34.210 42.510 ;
        RECT 35.410 41.240 35.550 43.900 ;
        RECT 36.330 41.240 36.470 43.900 ;
        RECT 37.550 42.910 37.690 45.570 ;
        RECT 38.460 42.910 38.600 45.570 ;
        RECT 39.820 45.480 40.330 45.790 ;
        RECT 39.820 44.210 39.960 45.480 ;
        RECT 41.160 44.210 41.300 46.310 ;
        RECT 42.080 44.210 42.220 46.310 ;
        RECT 43.300 45.880 43.440 47.980 ;
        RECT 44.210 45.880 44.350 47.980 ;
        RECT 45.570 47.890 46.080 48.200 ;
        RECT 45.570 46.620 45.710 47.890 ;
        RECT 46.910 46.620 47.050 49.330 ;
        RECT 47.830 46.620 47.970 50.590 ;
        RECT 49.050 48.290 49.190 50.590 ;
        RECT 49.960 49.750 50.100 50.590 ;
        RECT 51.180 50.340 51.580 50.740 ;
        RECT 49.960 49.330 50.350 49.750 ;
        RECT 51.320 49.720 51.460 50.340 ;
        RECT 52.660 49.750 52.800 50.590 ;
        RECT 51.230 49.400 51.550 49.720 ;
        RECT 49.960 48.290 50.100 49.330 ;
        RECT 48.960 47.980 49.280 48.290 ;
        RECT 49.870 47.980 50.190 48.290 ;
        RECT 51.320 48.200 51.460 49.400 ;
        RECT 52.400 49.330 52.800 49.750 ;
        RECT 45.180 46.310 45.710 46.620 ;
        RECT 46.820 46.310 47.140 46.620 ;
        RECT 47.730 46.310 48.050 46.620 ;
        RECT 43.210 45.570 43.530 45.880 ;
        RECT 44.120 45.570 44.440 45.880 ;
        RECT 45.570 45.790 45.710 46.310 ;
        RECT 39.430 43.900 39.960 44.210 ;
        RECT 41.070 43.900 41.390 44.210 ;
        RECT 41.980 43.900 42.300 44.210 ;
        RECT 37.460 42.600 37.780 42.910 ;
        RECT 38.370 42.600 38.690 42.910 ;
        RECT 39.820 42.820 39.960 43.900 ;
        RECT 33.680 40.930 34.210 41.240 ;
        RECT 35.320 40.930 35.640 41.240 ;
        RECT 36.230 40.930 36.550 41.240 ;
        RECT 31.710 40.190 32.030 40.500 ;
        RECT 32.620 40.190 32.940 40.500 ;
        RECT 34.070 40.410 34.210 40.930 ;
        RECT 27.930 38.520 28.460 38.830 ;
        RECT 29.570 38.520 29.890 38.830 ;
        RECT 30.480 38.520 30.800 38.830 ;
        RECT 25.960 37.780 26.280 38.090 ;
        RECT 26.870 37.780 27.190 38.090 ;
        RECT 28.320 38.000 28.460 38.520 ;
        RECT 22.180 36.110 22.710 36.420 ;
        RECT 23.820 36.110 24.140 36.420 ;
        RECT 24.730 36.110 25.050 36.420 ;
        RECT 20.210 35.370 20.530 35.680 ;
        RECT 21.120 35.370 21.440 35.680 ;
        RECT 22.570 35.590 22.710 36.110 ;
        RECT 16.430 33.700 16.960 34.010 ;
        RECT 18.070 33.700 18.390 34.010 ;
        RECT 18.980 33.700 19.300 34.010 ;
        RECT 14.460 32.960 14.780 33.270 ;
        RECT 15.370 32.960 15.690 33.270 ;
        RECT 16.820 33.180 16.960 33.700 ;
        RECT 10.680 31.290 11.210 31.600 ;
        RECT 12.320 31.290 12.640 31.600 ;
        RECT 13.230 31.290 13.550 31.600 ;
        RECT 8.710 30.550 9.030 30.860 ;
        RECT 9.620 30.550 9.940 30.860 ;
        RECT 11.070 30.770 11.210 31.290 ;
        RECT 4.930 28.880 5.460 29.190 ;
        RECT 6.570 28.880 6.890 29.190 ;
        RECT 7.480 28.880 7.800 29.190 ;
        RECT 2.960 27.740 3.280 28.050 ;
        RECT 3.870 27.740 4.190 28.050 ;
        RECT 5.320 27.960 5.460 28.880 ;
        RECT 1.280 25.700 1.540 26.020 ;
        RECT 1.350 23.610 1.500 25.700 ;
        RECT 3.050 25.640 3.190 27.740 ;
        RECT 3.960 25.640 4.100 27.740 ;
        RECT 5.320 27.650 5.830 27.960 ;
        RECT 5.320 26.380 5.460 27.650 ;
        RECT 6.660 26.380 6.800 28.880 ;
        RECT 7.580 26.380 7.720 28.880 ;
        RECT 8.800 28.050 8.940 30.550 ;
        RECT 9.710 28.050 9.850 30.550 ;
        RECT 11.070 30.460 11.580 30.770 ;
        RECT 11.070 29.190 11.210 30.460 ;
        RECT 12.410 29.190 12.550 31.290 ;
        RECT 13.330 29.190 13.470 31.290 ;
        RECT 14.550 30.860 14.690 32.960 ;
        RECT 15.460 30.860 15.600 32.960 ;
        RECT 16.820 32.870 17.330 33.180 ;
        RECT 16.820 31.600 16.960 32.870 ;
        RECT 18.160 31.600 18.300 33.700 ;
        RECT 19.080 31.600 19.220 33.700 ;
        RECT 20.300 33.270 20.440 35.370 ;
        RECT 21.210 33.270 21.350 35.370 ;
        RECT 22.570 35.280 23.080 35.590 ;
        RECT 22.570 34.010 22.710 35.280 ;
        RECT 23.910 34.010 24.050 36.110 ;
        RECT 24.830 34.010 24.970 36.110 ;
        RECT 26.050 35.680 26.190 37.780 ;
        RECT 26.960 35.680 27.100 37.780 ;
        RECT 28.320 37.690 28.830 38.000 ;
        RECT 28.320 36.420 28.460 37.690 ;
        RECT 29.660 36.420 29.800 38.520 ;
        RECT 30.580 36.420 30.720 38.520 ;
        RECT 31.800 38.090 31.940 40.190 ;
        RECT 32.710 38.090 32.850 40.190 ;
        RECT 34.070 40.100 34.580 40.410 ;
        RECT 34.070 38.830 34.210 40.100 ;
        RECT 35.410 38.830 35.550 40.930 ;
        RECT 36.330 38.830 36.470 40.930 ;
        RECT 37.550 40.500 37.690 42.600 ;
        RECT 38.460 40.500 38.600 42.600 ;
        RECT 39.820 42.510 40.330 42.820 ;
        RECT 39.820 41.240 39.960 42.510 ;
        RECT 41.160 41.240 41.300 43.900 ;
        RECT 42.080 41.240 42.220 43.900 ;
        RECT 43.300 42.910 43.440 45.570 ;
        RECT 44.210 42.910 44.350 45.570 ;
        RECT 45.570 45.480 46.080 45.790 ;
        RECT 45.570 44.210 45.710 45.480 ;
        RECT 46.910 44.210 47.050 46.310 ;
        RECT 47.830 44.210 47.970 46.310 ;
        RECT 49.050 45.880 49.190 47.980 ;
        RECT 49.960 45.880 50.100 47.980 ;
        RECT 51.320 47.890 51.830 48.200 ;
        RECT 51.320 46.620 51.460 47.890 ;
        RECT 52.660 46.620 52.800 49.330 ;
        RECT 53.580 46.620 53.720 50.590 ;
        RECT 54.800 48.290 54.940 50.590 ;
        RECT 55.710 49.750 55.850 50.590 ;
        RECT 56.940 50.340 57.340 50.740 ;
        RECT 55.710 49.330 56.100 49.750 ;
        RECT 57.070 49.720 57.210 50.340 ;
        RECT 58.410 49.750 58.550 50.590 ;
        RECT 56.980 49.400 57.300 49.720 ;
        RECT 55.710 48.290 55.850 49.330 ;
        RECT 54.710 47.980 55.030 48.290 ;
        RECT 55.620 47.980 55.940 48.290 ;
        RECT 57.070 48.200 57.210 49.400 ;
        RECT 58.150 49.330 58.550 49.750 ;
        RECT 50.930 46.310 51.460 46.620 ;
        RECT 52.570 46.310 52.890 46.620 ;
        RECT 53.480 46.310 53.800 46.620 ;
        RECT 48.960 45.570 49.280 45.880 ;
        RECT 49.870 45.570 50.190 45.880 ;
        RECT 51.320 45.790 51.460 46.310 ;
        RECT 45.180 43.900 45.710 44.210 ;
        RECT 46.820 43.900 47.140 44.210 ;
        RECT 47.730 43.900 48.050 44.210 ;
        RECT 43.210 42.600 43.530 42.910 ;
        RECT 44.120 42.600 44.440 42.910 ;
        RECT 45.570 42.820 45.710 43.900 ;
        RECT 39.430 40.930 39.960 41.240 ;
        RECT 41.070 40.930 41.390 41.240 ;
        RECT 41.980 40.930 42.300 41.240 ;
        RECT 37.460 40.190 37.780 40.500 ;
        RECT 38.370 40.190 38.690 40.500 ;
        RECT 39.820 40.410 39.960 40.930 ;
        RECT 33.680 38.520 34.210 38.830 ;
        RECT 35.320 38.520 35.640 38.830 ;
        RECT 36.230 38.520 36.550 38.830 ;
        RECT 31.710 37.780 32.030 38.090 ;
        RECT 32.620 37.780 32.940 38.090 ;
        RECT 34.070 38.000 34.210 38.520 ;
        RECT 27.930 36.110 28.460 36.420 ;
        RECT 29.570 36.110 29.890 36.420 ;
        RECT 30.480 36.110 30.800 36.420 ;
        RECT 25.960 35.370 26.280 35.680 ;
        RECT 26.870 35.370 27.190 35.680 ;
        RECT 28.320 35.590 28.460 36.110 ;
        RECT 22.180 33.700 22.710 34.010 ;
        RECT 23.820 33.700 24.140 34.010 ;
        RECT 24.730 33.700 25.050 34.010 ;
        RECT 20.210 32.960 20.530 33.270 ;
        RECT 21.120 32.960 21.440 33.270 ;
        RECT 22.570 33.180 22.710 33.700 ;
        RECT 16.430 31.290 16.960 31.600 ;
        RECT 18.070 31.290 18.390 31.600 ;
        RECT 18.980 31.290 19.300 31.600 ;
        RECT 14.460 30.550 14.780 30.860 ;
        RECT 15.370 30.550 15.690 30.860 ;
        RECT 16.820 30.770 16.960 31.290 ;
        RECT 10.680 28.880 11.210 29.190 ;
        RECT 12.320 28.880 12.640 29.190 ;
        RECT 13.230 28.880 13.550 29.190 ;
        RECT 8.710 27.740 9.030 28.050 ;
        RECT 9.620 27.740 9.940 28.050 ;
        RECT 11.070 27.960 11.210 28.880 ;
        RECT 4.930 26.070 5.460 26.380 ;
        RECT 6.570 26.070 6.890 26.380 ;
        RECT 7.480 26.070 7.800 26.380 ;
        RECT 2.960 25.330 3.280 25.640 ;
        RECT 3.870 25.330 4.190 25.640 ;
        RECT 5.320 25.550 5.460 26.070 ;
        RECT 1.290 23.290 1.550 23.610 ;
        RECT 1.350 21.200 1.500 23.290 ;
        RECT 3.050 23.230 3.190 25.330 ;
        RECT 3.960 23.230 4.100 25.330 ;
        RECT 5.320 25.240 5.830 25.550 ;
        RECT 5.320 23.970 5.460 25.240 ;
        RECT 6.660 23.970 6.800 26.070 ;
        RECT 7.580 23.970 7.720 26.070 ;
        RECT 8.800 25.640 8.940 27.740 ;
        RECT 9.710 25.640 9.850 27.740 ;
        RECT 11.070 27.650 11.580 27.960 ;
        RECT 11.070 26.380 11.210 27.650 ;
        RECT 12.410 26.380 12.550 28.880 ;
        RECT 13.330 26.380 13.470 28.880 ;
        RECT 14.550 28.050 14.690 30.550 ;
        RECT 15.460 28.050 15.600 30.550 ;
        RECT 16.820 30.460 17.330 30.770 ;
        RECT 16.820 29.190 16.960 30.460 ;
        RECT 18.160 29.190 18.300 31.290 ;
        RECT 19.080 29.190 19.220 31.290 ;
        RECT 20.300 30.860 20.440 32.960 ;
        RECT 21.210 30.860 21.350 32.960 ;
        RECT 22.570 32.870 23.080 33.180 ;
        RECT 22.570 31.600 22.710 32.870 ;
        RECT 23.910 31.600 24.050 33.700 ;
        RECT 24.830 31.600 24.970 33.700 ;
        RECT 26.050 33.270 26.190 35.370 ;
        RECT 26.960 33.270 27.100 35.370 ;
        RECT 28.320 35.280 28.830 35.590 ;
        RECT 28.320 34.010 28.460 35.280 ;
        RECT 29.660 34.010 29.800 36.110 ;
        RECT 30.580 34.010 30.720 36.110 ;
        RECT 31.800 35.680 31.940 37.780 ;
        RECT 32.710 35.680 32.850 37.780 ;
        RECT 34.070 37.690 34.580 38.000 ;
        RECT 34.070 36.420 34.210 37.690 ;
        RECT 35.410 36.420 35.550 38.520 ;
        RECT 36.330 36.420 36.470 38.520 ;
        RECT 37.550 38.090 37.690 40.190 ;
        RECT 38.460 38.090 38.600 40.190 ;
        RECT 39.820 40.100 40.330 40.410 ;
        RECT 39.820 38.830 39.960 40.100 ;
        RECT 41.160 38.830 41.300 40.930 ;
        RECT 42.080 38.830 42.220 40.930 ;
        RECT 43.300 40.500 43.440 42.600 ;
        RECT 44.210 40.500 44.350 42.600 ;
        RECT 45.570 42.510 46.080 42.820 ;
        RECT 45.570 41.240 45.710 42.510 ;
        RECT 46.910 41.240 47.050 43.900 ;
        RECT 47.830 41.240 47.970 43.900 ;
        RECT 49.050 42.910 49.190 45.570 ;
        RECT 49.960 42.910 50.100 45.570 ;
        RECT 51.320 45.480 51.830 45.790 ;
        RECT 51.320 44.210 51.460 45.480 ;
        RECT 52.660 44.210 52.800 46.310 ;
        RECT 53.580 44.210 53.720 46.310 ;
        RECT 54.800 45.880 54.940 47.980 ;
        RECT 55.710 45.880 55.850 47.980 ;
        RECT 57.070 47.890 57.580 48.200 ;
        RECT 57.070 46.620 57.210 47.890 ;
        RECT 58.410 46.620 58.550 49.330 ;
        RECT 59.330 46.620 59.470 50.590 ;
        RECT 60.550 48.290 60.690 50.590 ;
        RECT 61.460 49.750 61.600 50.590 ;
        RECT 62.690 50.330 63.090 50.730 ;
        RECT 61.460 49.330 61.850 49.750 ;
        RECT 62.820 49.720 62.960 50.330 ;
        RECT 64.160 49.750 64.300 50.590 ;
        RECT 62.730 49.400 63.050 49.720 ;
        RECT 61.460 48.290 61.600 49.330 ;
        RECT 60.460 47.980 60.780 48.290 ;
        RECT 61.370 47.980 61.690 48.290 ;
        RECT 62.820 48.200 62.960 49.400 ;
        RECT 63.900 49.330 64.300 49.750 ;
        RECT 56.680 46.310 57.210 46.620 ;
        RECT 58.320 46.310 58.640 46.620 ;
        RECT 59.230 46.310 59.550 46.620 ;
        RECT 54.710 45.570 55.030 45.880 ;
        RECT 55.620 45.570 55.940 45.880 ;
        RECT 57.070 45.790 57.210 46.310 ;
        RECT 50.930 43.900 51.460 44.210 ;
        RECT 52.570 43.900 52.890 44.210 ;
        RECT 53.480 43.900 53.800 44.210 ;
        RECT 48.960 42.600 49.280 42.910 ;
        RECT 49.870 42.600 50.190 42.910 ;
        RECT 51.320 42.820 51.460 43.900 ;
        RECT 45.180 40.930 45.710 41.240 ;
        RECT 46.820 40.930 47.140 41.240 ;
        RECT 47.730 40.930 48.050 41.240 ;
        RECT 43.210 40.190 43.530 40.500 ;
        RECT 44.120 40.190 44.440 40.500 ;
        RECT 45.570 40.410 45.710 40.930 ;
        RECT 39.430 38.520 39.960 38.830 ;
        RECT 41.070 38.520 41.390 38.830 ;
        RECT 41.980 38.520 42.300 38.830 ;
        RECT 37.460 37.780 37.780 38.090 ;
        RECT 38.370 37.780 38.690 38.090 ;
        RECT 39.820 38.000 39.960 38.520 ;
        RECT 33.680 36.110 34.210 36.420 ;
        RECT 35.320 36.110 35.640 36.420 ;
        RECT 36.230 36.110 36.550 36.420 ;
        RECT 31.710 35.370 32.030 35.680 ;
        RECT 32.620 35.370 32.940 35.680 ;
        RECT 34.070 35.590 34.210 36.110 ;
        RECT 27.930 33.700 28.460 34.010 ;
        RECT 29.570 33.700 29.890 34.010 ;
        RECT 30.480 33.700 30.800 34.010 ;
        RECT 25.960 32.960 26.280 33.270 ;
        RECT 26.870 32.960 27.190 33.270 ;
        RECT 28.320 33.180 28.460 33.700 ;
        RECT 22.180 31.290 22.710 31.600 ;
        RECT 23.820 31.290 24.140 31.600 ;
        RECT 24.730 31.290 25.050 31.600 ;
        RECT 20.210 30.550 20.530 30.860 ;
        RECT 21.120 30.550 21.440 30.860 ;
        RECT 22.570 30.770 22.710 31.290 ;
        RECT 16.430 28.880 16.960 29.190 ;
        RECT 18.070 28.880 18.390 29.190 ;
        RECT 18.980 28.880 19.300 29.190 ;
        RECT 14.460 27.740 14.780 28.050 ;
        RECT 15.370 27.740 15.690 28.050 ;
        RECT 16.820 27.960 16.960 28.880 ;
        RECT 10.680 26.070 11.210 26.380 ;
        RECT 12.320 26.070 12.640 26.380 ;
        RECT 13.230 26.070 13.550 26.380 ;
        RECT 8.710 25.330 9.030 25.640 ;
        RECT 9.620 25.330 9.940 25.640 ;
        RECT 11.070 25.550 11.210 26.070 ;
        RECT 4.930 23.660 5.460 23.970 ;
        RECT 6.570 23.660 6.890 23.970 ;
        RECT 7.480 23.660 7.800 23.970 ;
        RECT 2.960 22.920 3.280 23.230 ;
        RECT 3.870 22.920 4.190 23.230 ;
        RECT 5.320 23.140 5.460 23.660 ;
        RECT 1.290 20.880 1.550 21.200 ;
        RECT 1.350 18.790 1.500 20.880 ;
        RECT 3.050 20.820 3.190 22.920 ;
        RECT 3.960 20.820 4.100 22.920 ;
        RECT 5.320 22.830 5.830 23.140 ;
        RECT 5.320 21.560 5.460 22.830 ;
        RECT 6.660 21.560 6.800 23.660 ;
        RECT 7.580 21.560 7.720 23.660 ;
        RECT 8.800 23.230 8.940 25.330 ;
        RECT 9.710 23.230 9.850 25.330 ;
        RECT 11.070 25.240 11.580 25.550 ;
        RECT 11.070 23.970 11.210 25.240 ;
        RECT 12.410 23.970 12.550 26.070 ;
        RECT 13.330 23.970 13.470 26.070 ;
        RECT 14.550 25.640 14.690 27.740 ;
        RECT 15.460 25.640 15.600 27.740 ;
        RECT 16.820 27.650 17.330 27.960 ;
        RECT 16.820 26.380 16.960 27.650 ;
        RECT 18.160 26.380 18.300 28.880 ;
        RECT 19.080 26.380 19.220 28.880 ;
        RECT 20.300 28.050 20.440 30.550 ;
        RECT 21.210 28.050 21.350 30.550 ;
        RECT 22.570 30.460 23.080 30.770 ;
        RECT 22.570 29.190 22.710 30.460 ;
        RECT 23.910 29.190 24.050 31.290 ;
        RECT 24.830 29.190 24.970 31.290 ;
        RECT 26.050 30.860 26.190 32.960 ;
        RECT 26.960 30.860 27.100 32.960 ;
        RECT 28.320 32.870 28.830 33.180 ;
        RECT 28.320 31.600 28.460 32.870 ;
        RECT 29.660 31.600 29.800 33.700 ;
        RECT 30.580 31.600 30.720 33.700 ;
        RECT 31.800 33.270 31.940 35.370 ;
        RECT 32.710 33.270 32.850 35.370 ;
        RECT 34.070 35.280 34.580 35.590 ;
        RECT 34.070 34.010 34.210 35.280 ;
        RECT 35.410 34.010 35.550 36.110 ;
        RECT 36.330 34.010 36.470 36.110 ;
        RECT 37.550 35.680 37.690 37.780 ;
        RECT 38.460 35.680 38.600 37.780 ;
        RECT 39.820 37.690 40.330 38.000 ;
        RECT 39.820 36.420 39.960 37.690 ;
        RECT 41.160 36.420 41.300 38.520 ;
        RECT 42.080 36.420 42.220 38.520 ;
        RECT 43.300 38.090 43.440 40.190 ;
        RECT 44.210 38.090 44.350 40.190 ;
        RECT 45.570 40.100 46.080 40.410 ;
        RECT 45.570 38.830 45.710 40.100 ;
        RECT 46.910 38.830 47.050 40.930 ;
        RECT 47.830 38.830 47.970 40.930 ;
        RECT 49.050 40.500 49.190 42.600 ;
        RECT 49.960 40.500 50.100 42.600 ;
        RECT 51.320 42.510 51.830 42.820 ;
        RECT 51.320 41.240 51.460 42.510 ;
        RECT 52.660 41.240 52.800 43.900 ;
        RECT 53.580 41.240 53.720 43.900 ;
        RECT 54.800 42.910 54.940 45.570 ;
        RECT 55.710 42.910 55.850 45.570 ;
        RECT 57.070 45.480 57.580 45.790 ;
        RECT 57.070 44.210 57.210 45.480 ;
        RECT 58.410 44.210 58.550 46.310 ;
        RECT 59.330 44.210 59.470 46.310 ;
        RECT 60.550 45.880 60.690 47.980 ;
        RECT 61.460 45.880 61.600 47.980 ;
        RECT 62.820 47.890 63.330 48.200 ;
        RECT 62.820 46.620 62.960 47.890 ;
        RECT 64.160 46.620 64.300 49.330 ;
        RECT 65.080 46.620 65.220 50.590 ;
        RECT 66.300 48.290 66.440 50.590 ;
        RECT 67.210 49.750 67.350 50.590 ;
        RECT 68.430 50.340 68.830 50.740 ;
        RECT 67.210 49.330 67.600 49.750 ;
        RECT 68.570 49.720 68.710 50.340 ;
        RECT 69.910 49.750 70.050 50.590 ;
        RECT 68.480 49.400 68.800 49.720 ;
        RECT 67.210 48.290 67.350 49.330 ;
        RECT 66.210 47.980 66.530 48.290 ;
        RECT 67.120 47.980 67.440 48.290 ;
        RECT 68.570 48.200 68.710 49.400 ;
        RECT 69.650 49.330 70.050 49.750 ;
        RECT 62.430 46.310 62.960 46.620 ;
        RECT 64.070 46.310 64.390 46.620 ;
        RECT 64.980 46.310 65.300 46.620 ;
        RECT 60.460 45.570 60.780 45.880 ;
        RECT 61.370 45.570 61.690 45.880 ;
        RECT 62.820 45.790 62.960 46.310 ;
        RECT 56.680 43.900 57.210 44.210 ;
        RECT 58.320 43.900 58.640 44.210 ;
        RECT 59.230 43.900 59.550 44.210 ;
        RECT 54.710 42.600 55.030 42.910 ;
        RECT 55.620 42.600 55.940 42.910 ;
        RECT 57.070 42.820 57.210 43.900 ;
        RECT 50.930 40.930 51.460 41.240 ;
        RECT 52.570 40.930 52.890 41.240 ;
        RECT 53.480 40.930 53.800 41.240 ;
        RECT 48.960 40.190 49.280 40.500 ;
        RECT 49.870 40.190 50.190 40.500 ;
        RECT 51.320 40.410 51.460 40.930 ;
        RECT 45.180 38.520 45.710 38.830 ;
        RECT 46.820 38.520 47.140 38.830 ;
        RECT 47.730 38.520 48.050 38.830 ;
        RECT 43.210 37.780 43.530 38.090 ;
        RECT 44.120 37.780 44.440 38.090 ;
        RECT 45.570 38.000 45.710 38.520 ;
        RECT 39.430 36.110 39.960 36.420 ;
        RECT 41.070 36.110 41.390 36.420 ;
        RECT 41.980 36.110 42.300 36.420 ;
        RECT 37.460 35.370 37.780 35.680 ;
        RECT 38.370 35.370 38.690 35.680 ;
        RECT 39.820 35.590 39.960 36.110 ;
        RECT 33.680 33.700 34.210 34.010 ;
        RECT 35.320 33.700 35.640 34.010 ;
        RECT 36.230 33.700 36.550 34.010 ;
        RECT 31.710 32.960 32.030 33.270 ;
        RECT 32.620 32.960 32.940 33.270 ;
        RECT 34.070 33.180 34.210 33.700 ;
        RECT 27.930 31.290 28.460 31.600 ;
        RECT 29.570 31.290 29.890 31.600 ;
        RECT 30.480 31.290 30.800 31.600 ;
        RECT 25.960 30.550 26.280 30.860 ;
        RECT 26.870 30.550 27.190 30.860 ;
        RECT 28.320 30.770 28.460 31.290 ;
        RECT 22.180 28.880 22.710 29.190 ;
        RECT 23.820 28.880 24.140 29.190 ;
        RECT 24.730 28.880 25.050 29.190 ;
        RECT 20.210 27.740 20.530 28.050 ;
        RECT 21.120 27.740 21.440 28.050 ;
        RECT 22.570 27.960 22.710 28.880 ;
        RECT 16.430 26.070 16.960 26.380 ;
        RECT 18.070 26.070 18.390 26.380 ;
        RECT 18.980 26.070 19.300 26.380 ;
        RECT 14.460 25.330 14.780 25.640 ;
        RECT 15.370 25.330 15.690 25.640 ;
        RECT 16.820 25.550 16.960 26.070 ;
        RECT 10.680 23.660 11.210 23.970 ;
        RECT 12.320 23.660 12.640 23.970 ;
        RECT 13.230 23.660 13.550 23.970 ;
        RECT 8.710 22.920 9.030 23.230 ;
        RECT 9.620 22.920 9.940 23.230 ;
        RECT 11.070 23.140 11.210 23.660 ;
        RECT 4.930 21.250 5.460 21.560 ;
        RECT 6.570 21.250 6.890 21.560 ;
        RECT 7.480 21.250 7.800 21.560 ;
        RECT 2.960 20.510 3.280 20.820 ;
        RECT 3.870 20.510 4.190 20.820 ;
        RECT 5.320 20.730 5.460 21.250 ;
        RECT 1.290 18.470 1.550 18.790 ;
        RECT 1.350 16.380 1.500 18.470 ;
        RECT 3.050 18.410 3.190 20.510 ;
        RECT 3.960 18.410 4.100 20.510 ;
        RECT 5.320 20.420 5.830 20.730 ;
        RECT 5.320 19.150 5.460 20.420 ;
        RECT 6.660 19.150 6.800 21.250 ;
        RECT 7.580 19.150 7.720 21.250 ;
        RECT 8.800 20.820 8.940 22.920 ;
        RECT 9.710 20.820 9.850 22.920 ;
        RECT 11.070 22.830 11.580 23.140 ;
        RECT 11.070 21.560 11.210 22.830 ;
        RECT 12.410 21.560 12.550 23.660 ;
        RECT 13.330 21.560 13.470 23.660 ;
        RECT 14.550 23.230 14.690 25.330 ;
        RECT 15.460 23.230 15.600 25.330 ;
        RECT 16.820 25.240 17.330 25.550 ;
        RECT 16.820 23.970 16.960 25.240 ;
        RECT 18.160 23.970 18.300 26.070 ;
        RECT 19.080 23.970 19.220 26.070 ;
        RECT 20.300 25.640 20.440 27.740 ;
        RECT 21.210 25.640 21.350 27.740 ;
        RECT 22.570 27.650 23.080 27.960 ;
        RECT 22.570 26.380 22.710 27.650 ;
        RECT 23.910 26.380 24.050 28.880 ;
        RECT 24.830 26.380 24.970 28.880 ;
        RECT 26.050 28.050 26.190 30.550 ;
        RECT 26.960 28.050 27.100 30.550 ;
        RECT 28.320 30.460 28.830 30.770 ;
        RECT 28.320 29.190 28.460 30.460 ;
        RECT 29.660 29.190 29.800 31.290 ;
        RECT 30.580 29.190 30.720 31.290 ;
        RECT 31.800 30.860 31.940 32.960 ;
        RECT 32.710 30.860 32.850 32.960 ;
        RECT 34.070 32.870 34.580 33.180 ;
        RECT 34.070 31.600 34.210 32.870 ;
        RECT 35.410 31.600 35.550 33.700 ;
        RECT 36.330 31.600 36.470 33.700 ;
        RECT 37.550 33.270 37.690 35.370 ;
        RECT 38.460 33.270 38.600 35.370 ;
        RECT 39.820 35.280 40.330 35.590 ;
        RECT 39.820 34.010 39.960 35.280 ;
        RECT 41.160 34.010 41.300 36.110 ;
        RECT 42.080 34.010 42.220 36.110 ;
        RECT 43.300 35.680 43.440 37.780 ;
        RECT 44.210 35.680 44.350 37.780 ;
        RECT 45.570 37.690 46.080 38.000 ;
        RECT 45.570 36.420 45.710 37.690 ;
        RECT 46.910 36.420 47.050 38.520 ;
        RECT 47.830 36.420 47.970 38.520 ;
        RECT 49.050 38.090 49.190 40.190 ;
        RECT 49.960 38.090 50.100 40.190 ;
        RECT 51.320 40.100 51.830 40.410 ;
        RECT 51.320 38.830 51.460 40.100 ;
        RECT 52.660 38.830 52.800 40.930 ;
        RECT 53.580 38.830 53.720 40.930 ;
        RECT 54.800 40.500 54.940 42.600 ;
        RECT 55.710 40.500 55.850 42.600 ;
        RECT 57.070 42.510 57.580 42.820 ;
        RECT 57.070 41.240 57.210 42.510 ;
        RECT 58.410 41.240 58.550 43.900 ;
        RECT 59.330 41.240 59.470 43.900 ;
        RECT 60.550 42.910 60.690 45.570 ;
        RECT 61.460 42.910 61.600 45.570 ;
        RECT 62.820 45.480 63.330 45.790 ;
        RECT 62.820 44.210 62.960 45.480 ;
        RECT 64.160 44.210 64.300 46.310 ;
        RECT 65.080 44.210 65.220 46.310 ;
        RECT 66.300 45.880 66.440 47.980 ;
        RECT 67.210 45.880 67.350 47.980 ;
        RECT 68.570 47.890 69.080 48.200 ;
        RECT 68.570 46.620 68.710 47.890 ;
        RECT 69.910 46.620 70.050 49.330 ;
        RECT 70.830 46.620 70.970 50.590 ;
        RECT 72.050 48.290 72.190 50.590 ;
        RECT 72.960 49.750 73.100 50.590 ;
        RECT 74.180 50.340 74.580 50.740 ;
        RECT 72.960 49.330 73.350 49.750 ;
        RECT 74.320 49.720 74.460 50.340 ;
        RECT 75.660 49.750 75.800 50.590 ;
        RECT 74.230 49.400 74.550 49.720 ;
        RECT 72.960 48.290 73.100 49.330 ;
        RECT 71.960 47.980 72.280 48.290 ;
        RECT 72.870 47.980 73.190 48.290 ;
        RECT 74.320 48.200 74.460 49.400 ;
        RECT 75.400 49.330 75.800 49.750 ;
        RECT 68.180 46.310 68.710 46.620 ;
        RECT 69.820 46.310 70.140 46.620 ;
        RECT 70.730 46.310 71.050 46.620 ;
        RECT 66.210 45.570 66.530 45.880 ;
        RECT 67.120 45.570 67.440 45.880 ;
        RECT 68.570 45.790 68.710 46.310 ;
        RECT 62.430 43.900 62.960 44.210 ;
        RECT 64.070 43.900 64.390 44.210 ;
        RECT 64.980 43.900 65.300 44.210 ;
        RECT 60.460 42.600 60.780 42.910 ;
        RECT 61.370 42.600 61.690 42.910 ;
        RECT 62.820 42.820 62.960 43.900 ;
        RECT 56.680 40.930 57.210 41.240 ;
        RECT 58.320 40.930 58.640 41.240 ;
        RECT 59.230 40.930 59.550 41.240 ;
        RECT 54.710 40.190 55.030 40.500 ;
        RECT 55.620 40.190 55.940 40.500 ;
        RECT 57.070 40.410 57.210 40.930 ;
        RECT 50.930 38.520 51.460 38.830 ;
        RECT 52.570 38.520 52.890 38.830 ;
        RECT 53.480 38.520 53.800 38.830 ;
        RECT 48.960 37.780 49.280 38.090 ;
        RECT 49.870 37.780 50.190 38.090 ;
        RECT 51.320 38.000 51.460 38.520 ;
        RECT 45.180 36.110 45.710 36.420 ;
        RECT 46.820 36.110 47.140 36.420 ;
        RECT 47.730 36.110 48.050 36.420 ;
        RECT 43.210 35.370 43.530 35.680 ;
        RECT 44.120 35.370 44.440 35.680 ;
        RECT 45.570 35.590 45.710 36.110 ;
        RECT 39.430 33.700 39.960 34.010 ;
        RECT 41.070 33.700 41.390 34.010 ;
        RECT 41.980 33.700 42.300 34.010 ;
        RECT 37.460 32.960 37.780 33.270 ;
        RECT 38.370 32.960 38.690 33.270 ;
        RECT 39.820 33.180 39.960 33.700 ;
        RECT 33.680 31.290 34.210 31.600 ;
        RECT 35.320 31.290 35.640 31.600 ;
        RECT 36.230 31.290 36.550 31.600 ;
        RECT 31.710 30.550 32.030 30.860 ;
        RECT 32.620 30.550 32.940 30.860 ;
        RECT 34.070 30.770 34.210 31.290 ;
        RECT 27.930 28.880 28.460 29.190 ;
        RECT 29.570 28.880 29.890 29.190 ;
        RECT 30.480 28.880 30.800 29.190 ;
        RECT 25.960 27.740 26.280 28.050 ;
        RECT 26.870 27.740 27.190 28.050 ;
        RECT 28.320 27.960 28.460 28.880 ;
        RECT 22.180 26.070 22.710 26.380 ;
        RECT 23.820 26.070 24.140 26.380 ;
        RECT 24.730 26.070 25.050 26.380 ;
        RECT 20.210 25.330 20.530 25.640 ;
        RECT 21.120 25.330 21.440 25.640 ;
        RECT 22.570 25.550 22.710 26.070 ;
        RECT 16.430 23.660 16.960 23.970 ;
        RECT 18.070 23.660 18.390 23.970 ;
        RECT 18.980 23.660 19.300 23.970 ;
        RECT 14.460 22.920 14.780 23.230 ;
        RECT 15.370 22.920 15.690 23.230 ;
        RECT 16.820 23.140 16.960 23.660 ;
        RECT 10.680 21.250 11.210 21.560 ;
        RECT 12.320 21.250 12.640 21.560 ;
        RECT 13.230 21.250 13.550 21.560 ;
        RECT 8.710 20.510 9.030 20.820 ;
        RECT 9.620 20.510 9.940 20.820 ;
        RECT 11.070 20.730 11.210 21.250 ;
        RECT 4.930 18.840 5.460 19.150 ;
        RECT 6.570 18.840 6.890 19.150 ;
        RECT 7.480 18.840 7.800 19.150 ;
        RECT 2.960 18.100 3.280 18.410 ;
        RECT 3.870 18.100 4.190 18.410 ;
        RECT 5.320 18.320 5.460 18.840 ;
        RECT 1.290 16.060 1.550 16.380 ;
        RECT 1.350 13.970 1.500 16.060 ;
        RECT 3.050 16.000 3.190 18.100 ;
        RECT 3.960 16.000 4.100 18.100 ;
        RECT 5.320 18.010 5.830 18.320 ;
        RECT 5.320 16.740 5.460 18.010 ;
        RECT 6.660 16.740 6.800 18.840 ;
        RECT 7.580 16.740 7.720 18.840 ;
        RECT 8.800 18.410 8.940 20.510 ;
        RECT 9.710 18.410 9.850 20.510 ;
        RECT 11.070 20.420 11.580 20.730 ;
        RECT 11.070 19.150 11.210 20.420 ;
        RECT 12.410 19.150 12.550 21.250 ;
        RECT 13.330 19.150 13.470 21.250 ;
        RECT 14.550 20.820 14.690 22.920 ;
        RECT 15.460 20.820 15.600 22.920 ;
        RECT 16.820 22.830 17.330 23.140 ;
        RECT 16.820 21.560 16.960 22.830 ;
        RECT 18.160 21.560 18.300 23.660 ;
        RECT 19.080 21.560 19.220 23.660 ;
        RECT 20.300 23.230 20.440 25.330 ;
        RECT 21.210 23.230 21.350 25.330 ;
        RECT 22.570 25.240 23.080 25.550 ;
        RECT 22.570 23.970 22.710 25.240 ;
        RECT 23.910 23.970 24.050 26.070 ;
        RECT 24.830 23.970 24.970 26.070 ;
        RECT 26.050 25.640 26.190 27.740 ;
        RECT 26.960 25.640 27.100 27.740 ;
        RECT 28.320 27.650 28.830 27.960 ;
        RECT 28.320 26.380 28.460 27.650 ;
        RECT 29.660 26.380 29.800 28.880 ;
        RECT 30.580 26.380 30.720 28.880 ;
        RECT 31.800 28.050 31.940 30.550 ;
        RECT 32.710 28.050 32.850 30.550 ;
        RECT 34.070 30.460 34.580 30.770 ;
        RECT 34.070 29.190 34.210 30.460 ;
        RECT 35.410 29.190 35.550 31.290 ;
        RECT 36.330 29.190 36.470 31.290 ;
        RECT 37.550 30.860 37.690 32.960 ;
        RECT 38.460 30.860 38.600 32.960 ;
        RECT 39.820 32.870 40.330 33.180 ;
        RECT 39.820 31.600 39.960 32.870 ;
        RECT 41.160 31.600 41.300 33.700 ;
        RECT 42.080 31.600 42.220 33.700 ;
        RECT 43.300 33.270 43.440 35.370 ;
        RECT 44.210 33.270 44.350 35.370 ;
        RECT 45.570 35.280 46.080 35.590 ;
        RECT 45.570 34.010 45.710 35.280 ;
        RECT 46.910 34.010 47.050 36.110 ;
        RECT 47.830 34.010 47.970 36.110 ;
        RECT 49.050 35.680 49.190 37.780 ;
        RECT 49.960 35.680 50.100 37.780 ;
        RECT 51.320 37.690 51.830 38.000 ;
        RECT 51.320 36.420 51.460 37.690 ;
        RECT 52.660 36.420 52.800 38.520 ;
        RECT 53.580 36.420 53.720 38.520 ;
        RECT 54.800 38.090 54.940 40.190 ;
        RECT 55.710 38.090 55.850 40.190 ;
        RECT 57.070 40.100 57.580 40.410 ;
        RECT 57.070 38.830 57.210 40.100 ;
        RECT 58.410 38.830 58.550 40.930 ;
        RECT 59.330 38.830 59.470 40.930 ;
        RECT 60.550 40.500 60.690 42.600 ;
        RECT 61.460 40.500 61.600 42.600 ;
        RECT 62.820 42.510 63.330 42.820 ;
        RECT 62.820 41.240 62.960 42.510 ;
        RECT 64.160 41.240 64.300 43.900 ;
        RECT 65.080 41.240 65.220 43.900 ;
        RECT 66.300 42.910 66.440 45.570 ;
        RECT 67.210 42.910 67.350 45.570 ;
        RECT 68.570 45.480 69.080 45.790 ;
        RECT 68.570 44.210 68.710 45.480 ;
        RECT 69.910 44.210 70.050 46.310 ;
        RECT 70.830 44.210 70.970 46.310 ;
        RECT 72.050 45.880 72.190 47.980 ;
        RECT 72.960 45.880 73.100 47.980 ;
        RECT 74.320 47.890 74.830 48.200 ;
        RECT 74.320 46.620 74.460 47.890 ;
        RECT 75.660 46.620 75.800 49.330 ;
        RECT 76.580 46.620 76.720 50.590 ;
        RECT 77.800 48.290 77.940 50.590 ;
        RECT 78.710 49.750 78.850 50.590 ;
        RECT 79.930 50.340 80.330 50.740 ;
        RECT 78.710 49.330 79.100 49.750 ;
        RECT 80.070 49.720 80.210 50.340 ;
        RECT 81.410 49.750 81.550 50.590 ;
        RECT 79.980 49.400 80.300 49.720 ;
        RECT 78.710 48.290 78.850 49.330 ;
        RECT 77.710 47.980 78.030 48.290 ;
        RECT 78.620 47.980 78.940 48.290 ;
        RECT 80.070 48.200 80.210 49.400 ;
        RECT 81.150 49.330 81.550 49.750 ;
        RECT 73.930 46.310 74.460 46.620 ;
        RECT 75.570 46.310 75.890 46.620 ;
        RECT 76.480 46.310 76.800 46.620 ;
        RECT 71.960 45.570 72.280 45.880 ;
        RECT 72.870 45.570 73.190 45.880 ;
        RECT 74.320 45.790 74.460 46.310 ;
        RECT 68.180 43.900 68.710 44.210 ;
        RECT 69.820 43.900 70.140 44.210 ;
        RECT 70.730 43.900 71.050 44.210 ;
        RECT 66.210 42.600 66.530 42.910 ;
        RECT 67.120 42.600 67.440 42.910 ;
        RECT 68.570 42.820 68.710 43.900 ;
        RECT 62.430 40.930 62.960 41.240 ;
        RECT 64.070 40.930 64.390 41.240 ;
        RECT 64.980 40.930 65.300 41.240 ;
        RECT 60.460 40.190 60.780 40.500 ;
        RECT 61.370 40.190 61.690 40.500 ;
        RECT 62.820 40.410 62.960 40.930 ;
        RECT 56.680 38.520 57.210 38.830 ;
        RECT 58.320 38.520 58.640 38.830 ;
        RECT 59.230 38.520 59.550 38.830 ;
        RECT 54.710 37.780 55.030 38.090 ;
        RECT 55.620 37.780 55.940 38.090 ;
        RECT 57.070 38.000 57.210 38.520 ;
        RECT 50.930 36.110 51.460 36.420 ;
        RECT 52.570 36.110 52.890 36.420 ;
        RECT 53.480 36.110 53.800 36.420 ;
        RECT 48.960 35.370 49.280 35.680 ;
        RECT 49.870 35.370 50.190 35.680 ;
        RECT 51.320 35.590 51.460 36.110 ;
        RECT 45.180 33.700 45.710 34.010 ;
        RECT 46.820 33.700 47.140 34.010 ;
        RECT 47.730 33.700 48.050 34.010 ;
        RECT 43.210 32.960 43.530 33.270 ;
        RECT 44.120 32.960 44.440 33.270 ;
        RECT 45.570 33.180 45.710 33.700 ;
        RECT 39.430 31.290 39.960 31.600 ;
        RECT 41.070 31.290 41.390 31.600 ;
        RECT 41.980 31.290 42.300 31.600 ;
        RECT 37.460 30.550 37.780 30.860 ;
        RECT 38.370 30.550 38.690 30.860 ;
        RECT 39.820 30.770 39.960 31.290 ;
        RECT 33.680 28.880 34.210 29.190 ;
        RECT 35.320 28.880 35.640 29.190 ;
        RECT 36.230 28.880 36.550 29.190 ;
        RECT 31.710 27.740 32.030 28.050 ;
        RECT 32.620 27.740 32.940 28.050 ;
        RECT 34.070 27.960 34.210 28.880 ;
        RECT 27.930 26.070 28.460 26.380 ;
        RECT 29.570 26.070 29.890 26.380 ;
        RECT 30.480 26.070 30.800 26.380 ;
        RECT 25.960 25.330 26.280 25.640 ;
        RECT 26.870 25.330 27.190 25.640 ;
        RECT 28.320 25.550 28.460 26.070 ;
        RECT 22.180 23.660 22.710 23.970 ;
        RECT 23.820 23.660 24.140 23.970 ;
        RECT 24.730 23.660 25.050 23.970 ;
        RECT 20.210 22.920 20.530 23.230 ;
        RECT 21.120 22.920 21.440 23.230 ;
        RECT 22.570 23.140 22.710 23.660 ;
        RECT 16.430 21.250 16.960 21.560 ;
        RECT 18.070 21.250 18.390 21.560 ;
        RECT 18.980 21.250 19.300 21.560 ;
        RECT 14.460 20.510 14.780 20.820 ;
        RECT 15.370 20.510 15.690 20.820 ;
        RECT 16.820 20.730 16.960 21.250 ;
        RECT 10.680 18.840 11.210 19.150 ;
        RECT 12.320 18.840 12.640 19.150 ;
        RECT 13.230 18.840 13.550 19.150 ;
        RECT 8.710 18.100 9.030 18.410 ;
        RECT 9.620 18.100 9.940 18.410 ;
        RECT 11.070 18.320 11.210 18.840 ;
        RECT 4.930 16.430 5.460 16.740 ;
        RECT 6.570 16.430 6.890 16.740 ;
        RECT 7.480 16.430 7.800 16.740 ;
        RECT 2.960 15.690 3.280 16.000 ;
        RECT 3.870 15.690 4.190 16.000 ;
        RECT 5.320 15.910 5.460 16.430 ;
        RECT 1.290 13.650 1.550 13.970 ;
        RECT 1.350 11.560 1.500 13.650 ;
        RECT 3.050 13.590 3.190 15.690 ;
        RECT 3.960 13.590 4.100 15.690 ;
        RECT 5.320 15.600 5.830 15.910 ;
        RECT 5.320 14.330 5.460 15.600 ;
        RECT 6.660 14.330 6.800 16.430 ;
        RECT 7.580 14.330 7.720 16.430 ;
        RECT 8.800 16.000 8.940 18.100 ;
        RECT 9.710 16.000 9.850 18.100 ;
        RECT 11.070 18.010 11.580 18.320 ;
        RECT 11.070 16.740 11.210 18.010 ;
        RECT 12.410 16.740 12.550 18.840 ;
        RECT 13.330 16.740 13.470 18.840 ;
        RECT 14.550 18.410 14.690 20.510 ;
        RECT 15.460 18.410 15.600 20.510 ;
        RECT 16.820 20.420 17.330 20.730 ;
        RECT 16.820 19.150 16.960 20.420 ;
        RECT 18.160 19.150 18.300 21.250 ;
        RECT 19.080 19.150 19.220 21.250 ;
        RECT 20.300 20.820 20.440 22.920 ;
        RECT 21.210 20.820 21.350 22.920 ;
        RECT 22.570 22.830 23.080 23.140 ;
        RECT 22.570 21.560 22.710 22.830 ;
        RECT 23.910 21.560 24.050 23.660 ;
        RECT 24.830 21.560 24.970 23.660 ;
        RECT 26.050 23.230 26.190 25.330 ;
        RECT 26.960 23.230 27.100 25.330 ;
        RECT 28.320 25.240 28.830 25.550 ;
        RECT 28.320 23.970 28.460 25.240 ;
        RECT 29.660 23.970 29.800 26.070 ;
        RECT 30.580 23.970 30.720 26.070 ;
        RECT 31.800 25.640 31.940 27.740 ;
        RECT 32.710 25.640 32.850 27.740 ;
        RECT 34.070 27.650 34.580 27.960 ;
        RECT 34.070 26.380 34.210 27.650 ;
        RECT 35.410 26.380 35.550 28.880 ;
        RECT 36.330 26.380 36.470 28.880 ;
        RECT 37.550 28.050 37.690 30.550 ;
        RECT 38.460 28.050 38.600 30.550 ;
        RECT 39.820 30.460 40.330 30.770 ;
        RECT 39.820 29.190 39.960 30.460 ;
        RECT 41.160 29.190 41.300 31.290 ;
        RECT 42.080 29.190 42.220 31.290 ;
        RECT 43.300 30.860 43.440 32.960 ;
        RECT 44.210 30.860 44.350 32.960 ;
        RECT 45.570 32.870 46.080 33.180 ;
        RECT 45.570 31.600 45.710 32.870 ;
        RECT 46.910 31.600 47.050 33.700 ;
        RECT 47.830 31.600 47.970 33.700 ;
        RECT 49.050 33.270 49.190 35.370 ;
        RECT 49.960 33.270 50.100 35.370 ;
        RECT 51.320 35.280 51.830 35.590 ;
        RECT 51.320 34.010 51.460 35.280 ;
        RECT 52.660 34.010 52.800 36.110 ;
        RECT 53.580 34.010 53.720 36.110 ;
        RECT 54.800 35.680 54.940 37.780 ;
        RECT 55.710 35.680 55.850 37.780 ;
        RECT 57.070 37.690 57.580 38.000 ;
        RECT 57.070 36.420 57.210 37.690 ;
        RECT 58.410 36.420 58.550 38.520 ;
        RECT 59.330 36.420 59.470 38.520 ;
        RECT 60.550 38.090 60.690 40.190 ;
        RECT 61.460 38.090 61.600 40.190 ;
        RECT 62.820 40.100 63.330 40.410 ;
        RECT 62.820 38.830 62.960 40.100 ;
        RECT 64.160 38.830 64.300 40.930 ;
        RECT 65.080 38.830 65.220 40.930 ;
        RECT 66.300 40.500 66.440 42.600 ;
        RECT 67.210 40.500 67.350 42.600 ;
        RECT 68.570 42.510 69.080 42.820 ;
        RECT 68.570 41.240 68.710 42.510 ;
        RECT 69.910 41.240 70.050 43.900 ;
        RECT 70.830 41.240 70.970 43.900 ;
        RECT 72.050 42.910 72.190 45.570 ;
        RECT 72.960 42.910 73.100 45.570 ;
        RECT 74.320 45.480 74.830 45.790 ;
        RECT 74.320 44.210 74.460 45.480 ;
        RECT 75.660 44.210 75.800 46.310 ;
        RECT 76.580 44.210 76.720 46.310 ;
        RECT 77.800 45.880 77.940 47.980 ;
        RECT 78.710 45.880 78.850 47.980 ;
        RECT 80.070 47.890 80.580 48.200 ;
        RECT 80.070 46.620 80.210 47.890 ;
        RECT 81.410 46.620 81.550 49.330 ;
        RECT 82.330 46.620 82.470 50.590 ;
        RECT 83.550 48.290 83.690 50.590 ;
        RECT 84.460 49.750 84.600 50.590 ;
        RECT 85.670 50.340 86.070 50.740 ;
        RECT 84.460 49.330 84.850 49.750 ;
        RECT 85.820 49.720 85.960 50.340 ;
        RECT 87.160 49.750 87.300 50.590 ;
        RECT 85.730 49.400 86.050 49.720 ;
        RECT 84.460 48.290 84.600 49.330 ;
        RECT 83.460 47.980 83.780 48.290 ;
        RECT 84.370 47.980 84.690 48.290 ;
        RECT 85.820 48.200 85.960 49.400 ;
        RECT 86.900 49.330 87.300 49.750 ;
        RECT 79.680 46.310 80.210 46.620 ;
        RECT 81.320 46.310 81.640 46.620 ;
        RECT 82.230 46.310 82.550 46.620 ;
        RECT 77.710 45.570 78.030 45.880 ;
        RECT 78.620 45.570 78.940 45.880 ;
        RECT 80.070 45.790 80.210 46.310 ;
        RECT 73.930 43.900 74.460 44.210 ;
        RECT 75.570 43.900 75.890 44.210 ;
        RECT 76.480 43.900 76.800 44.210 ;
        RECT 71.960 42.600 72.280 42.910 ;
        RECT 72.870 42.600 73.190 42.910 ;
        RECT 74.320 42.820 74.460 43.900 ;
        RECT 68.180 40.930 68.710 41.240 ;
        RECT 69.820 40.930 70.140 41.240 ;
        RECT 70.730 40.930 71.050 41.240 ;
        RECT 66.210 40.190 66.530 40.500 ;
        RECT 67.120 40.190 67.440 40.500 ;
        RECT 68.570 40.410 68.710 40.930 ;
        RECT 62.430 38.520 62.960 38.830 ;
        RECT 64.070 38.520 64.390 38.830 ;
        RECT 64.980 38.520 65.300 38.830 ;
        RECT 60.460 37.780 60.780 38.090 ;
        RECT 61.370 37.780 61.690 38.090 ;
        RECT 62.820 38.000 62.960 38.520 ;
        RECT 56.680 36.110 57.210 36.420 ;
        RECT 58.320 36.110 58.640 36.420 ;
        RECT 59.230 36.110 59.550 36.420 ;
        RECT 54.710 35.370 55.030 35.680 ;
        RECT 55.620 35.370 55.940 35.680 ;
        RECT 57.070 35.590 57.210 36.110 ;
        RECT 50.930 33.700 51.460 34.010 ;
        RECT 52.570 33.700 52.890 34.010 ;
        RECT 53.480 33.700 53.800 34.010 ;
        RECT 48.960 32.960 49.280 33.270 ;
        RECT 49.870 32.960 50.190 33.270 ;
        RECT 51.320 33.180 51.460 33.700 ;
        RECT 45.180 31.290 45.710 31.600 ;
        RECT 46.820 31.290 47.140 31.600 ;
        RECT 47.730 31.290 48.050 31.600 ;
        RECT 43.210 30.550 43.530 30.860 ;
        RECT 44.120 30.550 44.440 30.860 ;
        RECT 45.570 30.770 45.710 31.290 ;
        RECT 39.430 28.880 39.960 29.190 ;
        RECT 41.070 28.880 41.390 29.190 ;
        RECT 41.980 28.880 42.300 29.190 ;
        RECT 37.460 27.740 37.780 28.050 ;
        RECT 38.370 27.740 38.690 28.050 ;
        RECT 39.820 27.960 39.960 28.880 ;
        RECT 33.680 26.070 34.210 26.380 ;
        RECT 35.320 26.070 35.640 26.380 ;
        RECT 36.230 26.070 36.550 26.380 ;
        RECT 31.710 25.330 32.030 25.640 ;
        RECT 32.620 25.330 32.940 25.640 ;
        RECT 34.070 25.550 34.210 26.070 ;
        RECT 27.930 23.660 28.460 23.970 ;
        RECT 29.570 23.660 29.890 23.970 ;
        RECT 30.480 23.660 30.800 23.970 ;
        RECT 25.960 22.920 26.280 23.230 ;
        RECT 26.870 22.920 27.190 23.230 ;
        RECT 28.320 23.140 28.460 23.660 ;
        RECT 22.180 21.250 22.710 21.560 ;
        RECT 23.820 21.250 24.140 21.560 ;
        RECT 24.730 21.250 25.050 21.560 ;
        RECT 20.210 20.510 20.530 20.820 ;
        RECT 21.120 20.510 21.440 20.820 ;
        RECT 22.570 20.730 22.710 21.250 ;
        RECT 16.430 18.840 16.960 19.150 ;
        RECT 18.070 18.840 18.390 19.150 ;
        RECT 18.980 18.840 19.300 19.150 ;
        RECT 14.460 18.100 14.780 18.410 ;
        RECT 15.370 18.100 15.690 18.410 ;
        RECT 16.820 18.320 16.960 18.840 ;
        RECT 10.680 16.430 11.210 16.740 ;
        RECT 12.320 16.430 12.640 16.740 ;
        RECT 13.230 16.430 13.550 16.740 ;
        RECT 8.710 15.690 9.030 16.000 ;
        RECT 9.620 15.690 9.940 16.000 ;
        RECT 11.070 15.910 11.210 16.430 ;
        RECT 4.930 14.020 5.460 14.330 ;
        RECT 6.570 14.020 6.890 14.330 ;
        RECT 7.480 14.020 7.800 14.330 ;
        RECT 2.960 13.280 3.280 13.590 ;
        RECT 3.870 13.280 4.190 13.590 ;
        RECT 5.320 13.500 5.460 14.020 ;
        RECT 1.280 11.240 1.540 11.560 ;
        RECT 1.350 9.150 1.500 11.240 ;
        RECT 3.050 11.180 3.190 13.280 ;
        RECT 3.960 11.180 4.100 13.280 ;
        RECT 5.320 13.190 5.830 13.500 ;
        RECT 5.320 11.920 5.460 13.190 ;
        RECT 6.660 11.920 6.800 14.020 ;
        RECT 7.580 11.920 7.720 14.020 ;
        RECT 8.800 13.590 8.940 15.690 ;
        RECT 9.710 13.590 9.850 15.690 ;
        RECT 11.070 15.600 11.580 15.910 ;
        RECT 11.070 14.330 11.210 15.600 ;
        RECT 12.410 14.330 12.550 16.430 ;
        RECT 13.330 14.330 13.470 16.430 ;
        RECT 14.550 16.000 14.690 18.100 ;
        RECT 15.460 16.000 15.600 18.100 ;
        RECT 16.820 18.010 17.330 18.320 ;
        RECT 16.820 16.740 16.960 18.010 ;
        RECT 18.160 16.740 18.300 18.840 ;
        RECT 19.080 16.740 19.220 18.840 ;
        RECT 20.300 18.410 20.440 20.510 ;
        RECT 21.210 18.410 21.350 20.510 ;
        RECT 22.570 20.420 23.080 20.730 ;
        RECT 22.570 19.150 22.710 20.420 ;
        RECT 23.910 19.150 24.050 21.250 ;
        RECT 24.830 19.150 24.970 21.250 ;
        RECT 26.050 20.820 26.190 22.920 ;
        RECT 26.960 20.820 27.100 22.920 ;
        RECT 28.320 22.830 28.830 23.140 ;
        RECT 28.320 21.560 28.460 22.830 ;
        RECT 29.660 21.560 29.800 23.660 ;
        RECT 30.580 21.560 30.720 23.660 ;
        RECT 31.800 23.230 31.940 25.330 ;
        RECT 32.710 23.230 32.850 25.330 ;
        RECT 34.070 25.240 34.580 25.550 ;
        RECT 34.070 23.970 34.210 25.240 ;
        RECT 35.410 23.970 35.550 26.070 ;
        RECT 36.330 23.970 36.470 26.070 ;
        RECT 37.550 25.640 37.690 27.740 ;
        RECT 38.460 25.640 38.600 27.740 ;
        RECT 39.820 27.650 40.330 27.960 ;
        RECT 39.820 26.380 39.960 27.650 ;
        RECT 41.160 26.380 41.300 28.880 ;
        RECT 42.080 26.380 42.220 28.880 ;
        RECT 43.300 28.050 43.440 30.550 ;
        RECT 44.210 28.050 44.350 30.550 ;
        RECT 45.570 30.460 46.080 30.770 ;
        RECT 45.570 29.190 45.710 30.460 ;
        RECT 46.910 29.190 47.050 31.290 ;
        RECT 47.830 29.190 47.970 31.290 ;
        RECT 49.050 30.860 49.190 32.960 ;
        RECT 49.960 30.860 50.100 32.960 ;
        RECT 51.320 32.870 51.830 33.180 ;
        RECT 51.320 31.600 51.460 32.870 ;
        RECT 52.660 31.600 52.800 33.700 ;
        RECT 53.580 31.600 53.720 33.700 ;
        RECT 54.800 33.270 54.940 35.370 ;
        RECT 55.710 33.270 55.850 35.370 ;
        RECT 57.070 35.280 57.580 35.590 ;
        RECT 57.070 34.010 57.210 35.280 ;
        RECT 58.410 34.010 58.550 36.110 ;
        RECT 59.330 34.010 59.470 36.110 ;
        RECT 60.550 35.680 60.690 37.780 ;
        RECT 61.460 35.680 61.600 37.780 ;
        RECT 62.820 37.690 63.330 38.000 ;
        RECT 62.820 36.420 62.960 37.690 ;
        RECT 64.160 36.420 64.300 38.520 ;
        RECT 65.080 36.420 65.220 38.520 ;
        RECT 66.300 38.090 66.440 40.190 ;
        RECT 67.210 38.090 67.350 40.190 ;
        RECT 68.570 40.100 69.080 40.410 ;
        RECT 68.570 38.830 68.710 40.100 ;
        RECT 69.910 38.830 70.050 40.930 ;
        RECT 70.830 38.830 70.970 40.930 ;
        RECT 72.050 40.500 72.190 42.600 ;
        RECT 72.960 40.500 73.100 42.600 ;
        RECT 74.320 42.510 74.830 42.820 ;
        RECT 74.320 41.240 74.460 42.510 ;
        RECT 75.660 41.240 75.800 43.900 ;
        RECT 76.580 41.240 76.720 43.900 ;
        RECT 77.800 42.910 77.940 45.570 ;
        RECT 78.710 42.910 78.850 45.570 ;
        RECT 80.070 45.480 80.580 45.790 ;
        RECT 80.070 44.210 80.210 45.480 ;
        RECT 81.410 44.210 81.550 46.310 ;
        RECT 82.330 44.210 82.470 46.310 ;
        RECT 83.550 45.880 83.690 47.980 ;
        RECT 84.460 45.880 84.600 47.980 ;
        RECT 85.820 47.890 86.330 48.200 ;
        RECT 85.820 46.620 85.960 47.890 ;
        RECT 87.160 46.620 87.300 49.330 ;
        RECT 88.080 46.620 88.220 50.590 ;
        RECT 89.300 48.290 89.440 50.590 ;
        RECT 90.210 49.750 90.350 50.590 ;
        RECT 91.420 50.340 91.820 50.740 ;
        RECT 90.210 49.330 90.600 49.750 ;
        RECT 91.570 49.720 91.710 50.340 ;
        RECT 92.910 49.750 93.050 50.590 ;
        RECT 91.480 49.400 91.800 49.720 ;
        RECT 90.210 48.290 90.350 49.330 ;
        RECT 89.210 47.980 89.530 48.290 ;
        RECT 90.120 47.980 90.440 48.290 ;
        RECT 91.570 48.200 91.710 49.400 ;
        RECT 92.650 49.330 93.050 49.750 ;
        RECT 85.430 46.310 85.960 46.620 ;
        RECT 87.070 46.310 87.390 46.620 ;
        RECT 87.980 46.310 88.300 46.620 ;
        RECT 83.460 45.570 83.780 45.880 ;
        RECT 84.370 45.570 84.690 45.880 ;
        RECT 85.820 45.790 85.960 46.310 ;
        RECT 79.680 43.900 80.210 44.210 ;
        RECT 81.320 43.900 81.640 44.210 ;
        RECT 82.230 43.900 82.550 44.210 ;
        RECT 77.710 42.600 78.030 42.910 ;
        RECT 78.620 42.600 78.940 42.910 ;
        RECT 80.070 42.820 80.210 43.900 ;
        RECT 73.930 40.930 74.460 41.240 ;
        RECT 75.570 40.930 75.890 41.240 ;
        RECT 76.480 40.930 76.800 41.240 ;
        RECT 71.960 40.190 72.280 40.500 ;
        RECT 72.870 40.190 73.190 40.500 ;
        RECT 74.320 40.410 74.460 40.930 ;
        RECT 68.180 38.520 68.710 38.830 ;
        RECT 69.820 38.520 70.140 38.830 ;
        RECT 70.730 38.520 71.050 38.830 ;
        RECT 66.210 37.780 66.530 38.090 ;
        RECT 67.120 37.780 67.440 38.090 ;
        RECT 68.570 38.000 68.710 38.520 ;
        RECT 62.430 36.110 62.960 36.420 ;
        RECT 64.070 36.110 64.390 36.420 ;
        RECT 64.980 36.110 65.300 36.420 ;
        RECT 60.460 35.370 60.780 35.680 ;
        RECT 61.370 35.370 61.690 35.680 ;
        RECT 62.820 35.590 62.960 36.110 ;
        RECT 56.680 33.700 57.210 34.010 ;
        RECT 58.320 33.700 58.640 34.010 ;
        RECT 59.230 33.700 59.550 34.010 ;
        RECT 54.710 32.960 55.030 33.270 ;
        RECT 55.620 32.960 55.940 33.270 ;
        RECT 57.070 33.180 57.210 33.700 ;
        RECT 50.930 31.290 51.460 31.600 ;
        RECT 52.570 31.290 52.890 31.600 ;
        RECT 53.480 31.290 53.800 31.600 ;
        RECT 48.960 30.550 49.280 30.860 ;
        RECT 49.870 30.550 50.190 30.860 ;
        RECT 51.320 30.770 51.460 31.290 ;
        RECT 45.180 28.880 45.710 29.190 ;
        RECT 46.820 28.880 47.140 29.190 ;
        RECT 47.730 28.880 48.050 29.190 ;
        RECT 43.210 27.740 43.530 28.050 ;
        RECT 44.120 27.740 44.440 28.050 ;
        RECT 45.570 27.960 45.710 28.880 ;
        RECT 39.430 26.070 39.960 26.380 ;
        RECT 41.070 26.070 41.390 26.380 ;
        RECT 41.980 26.070 42.300 26.380 ;
        RECT 37.460 25.330 37.780 25.640 ;
        RECT 38.370 25.330 38.690 25.640 ;
        RECT 39.820 25.550 39.960 26.070 ;
        RECT 33.680 23.660 34.210 23.970 ;
        RECT 35.320 23.660 35.640 23.970 ;
        RECT 36.230 23.660 36.550 23.970 ;
        RECT 31.710 22.920 32.030 23.230 ;
        RECT 32.620 22.920 32.940 23.230 ;
        RECT 34.070 23.140 34.210 23.660 ;
        RECT 27.930 21.250 28.460 21.560 ;
        RECT 29.570 21.250 29.890 21.560 ;
        RECT 30.480 21.250 30.800 21.560 ;
        RECT 25.960 20.510 26.280 20.820 ;
        RECT 26.870 20.510 27.190 20.820 ;
        RECT 28.320 20.730 28.460 21.250 ;
        RECT 22.180 18.840 22.710 19.150 ;
        RECT 23.820 18.840 24.140 19.150 ;
        RECT 24.730 18.840 25.050 19.150 ;
        RECT 20.210 18.100 20.530 18.410 ;
        RECT 21.120 18.100 21.440 18.410 ;
        RECT 22.570 18.320 22.710 18.840 ;
        RECT 16.430 16.430 16.960 16.740 ;
        RECT 18.070 16.430 18.390 16.740 ;
        RECT 18.980 16.430 19.300 16.740 ;
        RECT 14.460 15.690 14.780 16.000 ;
        RECT 15.370 15.690 15.690 16.000 ;
        RECT 16.820 15.910 16.960 16.430 ;
        RECT 10.680 14.020 11.210 14.330 ;
        RECT 12.320 14.020 12.640 14.330 ;
        RECT 13.230 14.020 13.550 14.330 ;
        RECT 8.710 13.280 9.030 13.590 ;
        RECT 9.620 13.280 9.940 13.590 ;
        RECT 11.070 13.500 11.210 14.020 ;
        RECT 4.930 11.610 5.460 11.920 ;
        RECT 6.570 11.610 6.890 11.920 ;
        RECT 7.480 11.610 7.800 11.920 ;
        RECT 2.960 10.870 3.280 11.180 ;
        RECT 3.870 10.870 4.190 11.180 ;
        RECT 5.320 11.090 5.460 11.610 ;
        RECT 1.290 8.830 1.550 9.150 ;
        RECT 1.350 6.330 1.500 8.830 ;
        RECT 3.050 8.360 3.190 10.870 ;
        RECT 3.960 8.360 4.100 10.870 ;
        RECT 5.320 10.780 5.830 11.090 ;
        RECT 5.320 9.510 5.460 10.780 ;
        RECT 6.660 9.510 6.800 11.610 ;
        RECT 7.580 9.510 7.720 11.610 ;
        RECT 8.800 11.180 8.940 13.280 ;
        RECT 9.710 11.180 9.850 13.280 ;
        RECT 11.070 13.190 11.580 13.500 ;
        RECT 11.070 11.920 11.210 13.190 ;
        RECT 12.410 11.920 12.550 14.020 ;
        RECT 13.330 11.920 13.470 14.020 ;
        RECT 14.550 13.590 14.690 15.690 ;
        RECT 15.460 13.590 15.600 15.690 ;
        RECT 16.820 15.600 17.330 15.910 ;
        RECT 16.820 14.330 16.960 15.600 ;
        RECT 18.160 14.330 18.300 16.430 ;
        RECT 19.080 14.330 19.220 16.430 ;
        RECT 20.300 16.000 20.440 18.100 ;
        RECT 21.210 16.000 21.350 18.100 ;
        RECT 22.570 18.010 23.080 18.320 ;
        RECT 22.570 16.740 22.710 18.010 ;
        RECT 23.910 16.740 24.050 18.840 ;
        RECT 24.830 16.740 24.970 18.840 ;
        RECT 26.050 18.410 26.190 20.510 ;
        RECT 26.960 18.410 27.100 20.510 ;
        RECT 28.320 20.420 28.830 20.730 ;
        RECT 28.320 19.150 28.460 20.420 ;
        RECT 29.660 19.150 29.800 21.250 ;
        RECT 30.580 19.150 30.720 21.250 ;
        RECT 31.800 20.820 31.940 22.920 ;
        RECT 32.710 20.820 32.850 22.920 ;
        RECT 34.070 22.830 34.580 23.140 ;
        RECT 34.070 21.560 34.210 22.830 ;
        RECT 35.410 21.560 35.550 23.660 ;
        RECT 36.330 21.560 36.470 23.660 ;
        RECT 37.550 23.230 37.690 25.330 ;
        RECT 38.460 23.230 38.600 25.330 ;
        RECT 39.820 25.240 40.330 25.550 ;
        RECT 39.820 23.970 39.960 25.240 ;
        RECT 41.160 23.970 41.300 26.070 ;
        RECT 42.080 23.970 42.220 26.070 ;
        RECT 43.300 25.640 43.440 27.740 ;
        RECT 44.210 25.640 44.350 27.740 ;
        RECT 45.570 27.650 46.080 27.960 ;
        RECT 45.570 26.380 45.710 27.650 ;
        RECT 46.910 26.380 47.050 28.880 ;
        RECT 47.830 26.380 47.970 28.880 ;
        RECT 49.050 28.050 49.190 30.550 ;
        RECT 49.960 28.050 50.100 30.550 ;
        RECT 51.320 30.460 51.830 30.770 ;
        RECT 51.320 29.190 51.460 30.460 ;
        RECT 52.660 29.190 52.800 31.290 ;
        RECT 53.580 29.190 53.720 31.290 ;
        RECT 54.800 30.860 54.940 32.960 ;
        RECT 55.710 30.860 55.850 32.960 ;
        RECT 57.070 32.870 57.580 33.180 ;
        RECT 57.070 31.600 57.210 32.870 ;
        RECT 58.410 31.600 58.550 33.700 ;
        RECT 59.330 31.600 59.470 33.700 ;
        RECT 60.550 33.270 60.690 35.370 ;
        RECT 61.460 33.270 61.600 35.370 ;
        RECT 62.820 35.280 63.330 35.590 ;
        RECT 62.820 34.010 62.960 35.280 ;
        RECT 64.160 34.010 64.300 36.110 ;
        RECT 65.080 34.010 65.220 36.110 ;
        RECT 66.300 35.680 66.440 37.780 ;
        RECT 67.210 35.680 67.350 37.780 ;
        RECT 68.570 37.690 69.080 38.000 ;
        RECT 68.570 36.420 68.710 37.690 ;
        RECT 69.910 36.420 70.050 38.520 ;
        RECT 70.830 36.420 70.970 38.520 ;
        RECT 72.050 38.090 72.190 40.190 ;
        RECT 72.960 38.090 73.100 40.190 ;
        RECT 74.320 40.100 74.830 40.410 ;
        RECT 74.320 38.830 74.460 40.100 ;
        RECT 75.660 38.830 75.800 40.930 ;
        RECT 76.580 38.830 76.720 40.930 ;
        RECT 77.800 40.500 77.940 42.600 ;
        RECT 78.710 40.500 78.850 42.600 ;
        RECT 80.070 42.510 80.580 42.820 ;
        RECT 80.070 41.240 80.210 42.510 ;
        RECT 81.410 41.240 81.550 43.900 ;
        RECT 82.330 41.240 82.470 43.900 ;
        RECT 83.550 42.910 83.690 45.570 ;
        RECT 84.460 42.910 84.600 45.570 ;
        RECT 85.820 45.480 86.330 45.790 ;
        RECT 85.820 44.210 85.960 45.480 ;
        RECT 87.160 44.210 87.300 46.310 ;
        RECT 88.080 44.210 88.220 46.310 ;
        RECT 89.300 45.880 89.440 47.980 ;
        RECT 90.210 45.880 90.350 47.980 ;
        RECT 91.570 47.890 92.080 48.200 ;
        RECT 91.570 46.620 91.710 47.890 ;
        RECT 92.910 46.620 93.050 49.330 ;
        RECT 93.830 46.620 93.970 50.590 ;
        RECT 91.180 46.310 91.710 46.620 ;
        RECT 92.820 46.310 93.140 46.620 ;
        RECT 93.730 46.310 94.050 46.620 ;
        RECT 89.210 45.570 89.530 45.880 ;
        RECT 90.120 45.570 90.440 45.880 ;
        RECT 91.570 45.790 91.710 46.310 ;
        RECT 85.430 43.900 85.960 44.210 ;
        RECT 87.070 43.900 87.390 44.210 ;
        RECT 87.980 43.900 88.300 44.210 ;
        RECT 83.460 42.600 83.780 42.910 ;
        RECT 84.370 42.600 84.690 42.910 ;
        RECT 85.820 42.820 85.960 43.900 ;
        RECT 79.680 40.930 80.210 41.240 ;
        RECT 81.320 40.930 81.640 41.240 ;
        RECT 82.230 40.930 82.550 41.240 ;
        RECT 77.710 40.190 78.030 40.500 ;
        RECT 78.620 40.190 78.940 40.500 ;
        RECT 80.070 40.410 80.210 40.930 ;
        RECT 73.930 38.520 74.460 38.830 ;
        RECT 75.570 38.520 75.890 38.830 ;
        RECT 76.480 38.520 76.800 38.830 ;
        RECT 71.960 37.780 72.280 38.090 ;
        RECT 72.870 37.780 73.190 38.090 ;
        RECT 74.320 38.000 74.460 38.520 ;
        RECT 68.180 36.110 68.710 36.420 ;
        RECT 69.820 36.110 70.140 36.420 ;
        RECT 70.730 36.110 71.050 36.420 ;
        RECT 66.210 35.370 66.530 35.680 ;
        RECT 67.120 35.370 67.440 35.680 ;
        RECT 68.570 35.590 68.710 36.110 ;
        RECT 62.430 33.700 62.960 34.010 ;
        RECT 64.070 33.700 64.390 34.010 ;
        RECT 64.980 33.700 65.300 34.010 ;
        RECT 60.460 32.960 60.780 33.270 ;
        RECT 61.370 32.960 61.690 33.270 ;
        RECT 62.820 33.180 62.960 33.700 ;
        RECT 56.680 31.290 57.210 31.600 ;
        RECT 58.320 31.290 58.640 31.600 ;
        RECT 59.230 31.290 59.550 31.600 ;
        RECT 54.710 30.550 55.030 30.860 ;
        RECT 55.620 30.550 55.940 30.860 ;
        RECT 57.070 30.770 57.210 31.290 ;
        RECT 50.930 28.880 51.460 29.190 ;
        RECT 52.570 28.880 52.890 29.190 ;
        RECT 53.480 28.880 53.800 29.190 ;
        RECT 48.960 27.740 49.280 28.050 ;
        RECT 49.870 27.740 50.190 28.050 ;
        RECT 51.320 27.960 51.460 28.880 ;
        RECT 45.180 26.070 45.710 26.380 ;
        RECT 46.820 26.070 47.140 26.380 ;
        RECT 47.730 26.070 48.050 26.380 ;
        RECT 43.210 25.330 43.530 25.640 ;
        RECT 44.120 25.330 44.440 25.640 ;
        RECT 45.570 25.550 45.710 26.070 ;
        RECT 39.430 23.660 39.960 23.970 ;
        RECT 41.070 23.660 41.390 23.970 ;
        RECT 41.980 23.660 42.300 23.970 ;
        RECT 37.460 22.920 37.780 23.230 ;
        RECT 38.370 22.920 38.690 23.230 ;
        RECT 39.820 23.140 39.960 23.660 ;
        RECT 33.680 21.250 34.210 21.560 ;
        RECT 35.320 21.250 35.640 21.560 ;
        RECT 36.230 21.250 36.550 21.560 ;
        RECT 31.710 20.510 32.030 20.820 ;
        RECT 32.620 20.510 32.940 20.820 ;
        RECT 34.070 20.730 34.210 21.250 ;
        RECT 27.930 18.840 28.460 19.150 ;
        RECT 29.570 18.840 29.890 19.150 ;
        RECT 30.480 18.840 30.800 19.150 ;
        RECT 25.960 18.100 26.280 18.410 ;
        RECT 26.870 18.100 27.190 18.410 ;
        RECT 28.320 18.320 28.460 18.840 ;
        RECT 22.180 16.430 22.710 16.740 ;
        RECT 23.820 16.430 24.140 16.740 ;
        RECT 24.730 16.430 25.050 16.740 ;
        RECT 20.210 15.690 20.530 16.000 ;
        RECT 21.120 15.690 21.440 16.000 ;
        RECT 22.570 15.910 22.710 16.430 ;
        RECT 16.430 14.020 16.960 14.330 ;
        RECT 18.070 14.020 18.390 14.330 ;
        RECT 18.980 14.020 19.300 14.330 ;
        RECT 14.460 13.280 14.780 13.590 ;
        RECT 15.370 13.280 15.690 13.590 ;
        RECT 16.820 13.500 16.960 14.020 ;
        RECT 10.680 11.610 11.210 11.920 ;
        RECT 12.320 11.610 12.640 11.920 ;
        RECT 13.230 11.610 13.550 11.920 ;
        RECT 8.710 10.870 9.030 11.180 ;
        RECT 9.620 10.870 9.940 11.180 ;
        RECT 11.070 11.090 11.210 11.610 ;
        RECT 4.930 9.200 5.460 9.510 ;
        RECT 6.570 9.200 6.890 9.510 ;
        RECT 7.480 9.200 7.800 9.510 ;
        RECT 2.960 8.050 3.280 8.360 ;
        RECT 3.870 8.050 4.190 8.360 ;
        RECT 5.320 8.270 5.460 9.200 ;
        RECT 1.280 6.010 1.540 6.330 ;
        RECT 1.350 3.920 1.500 6.010 ;
        RECT 3.050 5.950 3.190 8.050 ;
        RECT 3.960 5.950 4.100 8.050 ;
        RECT 5.320 7.960 5.830 8.270 ;
        RECT 5.320 6.690 5.460 7.960 ;
        RECT 6.660 6.690 6.800 9.200 ;
        RECT 7.580 6.690 7.720 9.200 ;
        RECT 8.800 8.360 8.940 10.870 ;
        RECT 9.710 8.360 9.850 10.870 ;
        RECT 11.070 10.780 11.580 11.090 ;
        RECT 11.070 9.510 11.210 10.780 ;
        RECT 12.410 9.510 12.550 11.610 ;
        RECT 13.330 9.510 13.470 11.610 ;
        RECT 14.550 11.180 14.690 13.280 ;
        RECT 15.460 11.180 15.600 13.280 ;
        RECT 16.820 13.190 17.330 13.500 ;
        RECT 16.820 11.920 16.960 13.190 ;
        RECT 18.160 11.920 18.300 14.020 ;
        RECT 19.080 11.920 19.220 14.020 ;
        RECT 20.300 13.590 20.440 15.690 ;
        RECT 21.210 13.590 21.350 15.690 ;
        RECT 22.570 15.600 23.080 15.910 ;
        RECT 22.570 14.330 22.710 15.600 ;
        RECT 23.910 14.330 24.050 16.430 ;
        RECT 24.830 14.330 24.970 16.430 ;
        RECT 26.050 16.000 26.190 18.100 ;
        RECT 26.960 16.000 27.100 18.100 ;
        RECT 28.320 18.010 28.830 18.320 ;
        RECT 28.320 16.740 28.460 18.010 ;
        RECT 29.660 16.740 29.800 18.840 ;
        RECT 30.580 16.740 30.720 18.840 ;
        RECT 31.800 18.410 31.940 20.510 ;
        RECT 32.710 18.410 32.850 20.510 ;
        RECT 34.070 20.420 34.580 20.730 ;
        RECT 34.070 19.150 34.210 20.420 ;
        RECT 35.410 19.150 35.550 21.250 ;
        RECT 36.330 19.150 36.470 21.250 ;
        RECT 37.550 20.820 37.690 22.920 ;
        RECT 38.460 20.820 38.600 22.920 ;
        RECT 39.820 22.830 40.330 23.140 ;
        RECT 39.820 21.560 39.960 22.830 ;
        RECT 41.160 21.560 41.300 23.660 ;
        RECT 42.080 21.560 42.220 23.660 ;
        RECT 43.300 23.230 43.440 25.330 ;
        RECT 44.210 23.230 44.350 25.330 ;
        RECT 45.570 25.240 46.080 25.550 ;
        RECT 45.570 23.970 45.710 25.240 ;
        RECT 46.910 23.970 47.050 26.070 ;
        RECT 47.830 23.970 47.970 26.070 ;
        RECT 49.050 25.640 49.190 27.740 ;
        RECT 49.960 25.640 50.100 27.740 ;
        RECT 51.320 27.650 51.830 27.960 ;
        RECT 51.320 26.380 51.460 27.650 ;
        RECT 52.660 26.380 52.800 28.880 ;
        RECT 53.580 26.380 53.720 28.880 ;
        RECT 54.800 28.050 54.940 30.550 ;
        RECT 55.710 28.050 55.850 30.550 ;
        RECT 57.070 30.460 57.580 30.770 ;
        RECT 57.070 29.190 57.210 30.460 ;
        RECT 58.410 29.190 58.550 31.290 ;
        RECT 59.330 29.190 59.470 31.290 ;
        RECT 60.550 30.860 60.690 32.960 ;
        RECT 61.460 30.860 61.600 32.960 ;
        RECT 62.820 32.870 63.330 33.180 ;
        RECT 62.820 31.600 62.960 32.870 ;
        RECT 64.160 31.600 64.300 33.700 ;
        RECT 65.080 31.600 65.220 33.700 ;
        RECT 66.300 33.270 66.440 35.370 ;
        RECT 67.210 33.270 67.350 35.370 ;
        RECT 68.570 35.280 69.080 35.590 ;
        RECT 68.570 34.010 68.710 35.280 ;
        RECT 69.910 34.010 70.050 36.110 ;
        RECT 70.830 34.010 70.970 36.110 ;
        RECT 72.050 35.680 72.190 37.780 ;
        RECT 72.960 35.680 73.100 37.780 ;
        RECT 74.320 37.690 74.830 38.000 ;
        RECT 74.320 36.420 74.460 37.690 ;
        RECT 75.660 36.420 75.800 38.520 ;
        RECT 76.580 36.420 76.720 38.520 ;
        RECT 77.800 38.090 77.940 40.190 ;
        RECT 78.710 38.090 78.850 40.190 ;
        RECT 80.070 40.100 80.580 40.410 ;
        RECT 80.070 38.830 80.210 40.100 ;
        RECT 81.410 38.830 81.550 40.930 ;
        RECT 82.330 38.830 82.470 40.930 ;
        RECT 83.550 40.500 83.690 42.600 ;
        RECT 84.460 40.500 84.600 42.600 ;
        RECT 85.820 42.510 86.330 42.820 ;
        RECT 85.820 41.240 85.960 42.510 ;
        RECT 87.160 41.240 87.300 43.900 ;
        RECT 88.080 41.240 88.220 43.900 ;
        RECT 89.300 42.910 89.440 45.570 ;
        RECT 90.210 42.910 90.350 45.570 ;
        RECT 91.570 45.480 92.080 45.790 ;
        RECT 91.570 44.210 91.710 45.480 ;
        RECT 92.910 44.210 93.050 46.310 ;
        RECT 93.830 44.210 93.970 46.310 ;
        RECT 91.180 43.900 91.710 44.210 ;
        RECT 92.820 43.900 93.140 44.210 ;
        RECT 93.730 43.900 94.050 44.210 ;
        RECT 89.210 42.600 89.530 42.910 ;
        RECT 90.120 42.600 90.440 42.910 ;
        RECT 91.570 42.820 91.710 43.900 ;
        RECT 85.430 40.930 85.960 41.240 ;
        RECT 87.070 40.930 87.390 41.240 ;
        RECT 87.980 40.930 88.300 41.240 ;
        RECT 83.460 40.190 83.780 40.500 ;
        RECT 84.370 40.190 84.690 40.500 ;
        RECT 85.820 40.410 85.960 40.930 ;
        RECT 79.680 38.520 80.210 38.830 ;
        RECT 81.320 38.520 81.640 38.830 ;
        RECT 82.230 38.520 82.550 38.830 ;
        RECT 77.710 37.780 78.030 38.090 ;
        RECT 78.620 37.780 78.940 38.090 ;
        RECT 80.070 38.000 80.210 38.520 ;
        RECT 73.930 36.110 74.460 36.420 ;
        RECT 75.570 36.110 75.890 36.420 ;
        RECT 76.480 36.110 76.800 36.420 ;
        RECT 71.960 35.370 72.280 35.680 ;
        RECT 72.870 35.370 73.190 35.680 ;
        RECT 74.320 35.590 74.460 36.110 ;
        RECT 68.180 33.700 68.710 34.010 ;
        RECT 69.820 33.700 70.140 34.010 ;
        RECT 70.730 33.700 71.050 34.010 ;
        RECT 66.210 32.960 66.530 33.270 ;
        RECT 67.120 32.960 67.440 33.270 ;
        RECT 68.570 33.180 68.710 33.700 ;
        RECT 62.430 31.290 62.960 31.600 ;
        RECT 64.070 31.290 64.390 31.600 ;
        RECT 64.980 31.290 65.300 31.600 ;
        RECT 60.460 30.550 60.780 30.860 ;
        RECT 61.370 30.550 61.690 30.860 ;
        RECT 62.820 30.770 62.960 31.290 ;
        RECT 56.680 28.880 57.210 29.190 ;
        RECT 58.320 28.880 58.640 29.190 ;
        RECT 59.230 28.880 59.550 29.190 ;
        RECT 54.710 27.740 55.030 28.050 ;
        RECT 55.620 27.740 55.940 28.050 ;
        RECT 57.070 27.960 57.210 28.880 ;
        RECT 50.930 26.070 51.460 26.380 ;
        RECT 52.570 26.070 52.890 26.380 ;
        RECT 53.480 26.070 53.800 26.380 ;
        RECT 48.960 25.330 49.280 25.640 ;
        RECT 49.870 25.330 50.190 25.640 ;
        RECT 51.320 25.550 51.460 26.070 ;
        RECT 45.180 23.660 45.710 23.970 ;
        RECT 46.820 23.660 47.140 23.970 ;
        RECT 47.730 23.660 48.050 23.970 ;
        RECT 43.210 22.920 43.530 23.230 ;
        RECT 44.120 22.920 44.440 23.230 ;
        RECT 45.570 23.140 45.710 23.660 ;
        RECT 39.430 21.250 39.960 21.560 ;
        RECT 41.070 21.250 41.390 21.560 ;
        RECT 41.980 21.250 42.300 21.560 ;
        RECT 37.460 20.510 37.780 20.820 ;
        RECT 38.370 20.510 38.690 20.820 ;
        RECT 39.820 20.730 39.960 21.250 ;
        RECT 33.680 18.840 34.210 19.150 ;
        RECT 35.320 18.840 35.640 19.150 ;
        RECT 36.230 18.840 36.550 19.150 ;
        RECT 31.710 18.100 32.030 18.410 ;
        RECT 32.620 18.100 32.940 18.410 ;
        RECT 34.070 18.320 34.210 18.840 ;
        RECT 27.930 16.430 28.460 16.740 ;
        RECT 29.570 16.430 29.890 16.740 ;
        RECT 30.480 16.430 30.800 16.740 ;
        RECT 25.960 15.690 26.280 16.000 ;
        RECT 26.870 15.690 27.190 16.000 ;
        RECT 28.320 15.910 28.460 16.430 ;
        RECT 22.180 14.020 22.710 14.330 ;
        RECT 23.820 14.020 24.140 14.330 ;
        RECT 24.730 14.020 25.050 14.330 ;
        RECT 20.210 13.280 20.530 13.590 ;
        RECT 21.120 13.280 21.440 13.590 ;
        RECT 22.570 13.500 22.710 14.020 ;
        RECT 16.430 11.610 16.960 11.920 ;
        RECT 18.070 11.610 18.390 11.920 ;
        RECT 18.980 11.610 19.300 11.920 ;
        RECT 14.460 10.870 14.780 11.180 ;
        RECT 15.370 10.870 15.690 11.180 ;
        RECT 16.820 11.090 16.960 11.610 ;
        RECT 10.680 9.200 11.210 9.510 ;
        RECT 12.320 9.200 12.640 9.510 ;
        RECT 13.230 9.200 13.550 9.510 ;
        RECT 8.710 8.050 9.030 8.360 ;
        RECT 9.620 8.050 9.940 8.360 ;
        RECT 11.070 8.270 11.210 9.200 ;
        RECT 4.930 6.380 5.460 6.690 ;
        RECT 6.570 6.380 6.890 6.690 ;
        RECT 7.480 6.380 7.800 6.690 ;
        RECT 2.960 5.640 3.280 5.950 ;
        RECT 3.870 5.640 4.190 5.950 ;
        RECT 5.320 5.860 5.460 6.380 ;
        RECT 1.300 3.600 1.560 3.920 ;
        RECT 1.350 1.510 1.500 3.600 ;
        RECT 3.050 3.540 3.190 5.640 ;
        RECT 3.960 3.540 4.100 5.640 ;
        RECT 5.320 5.550 5.830 5.860 ;
        RECT 5.320 4.280 5.460 5.550 ;
        RECT 6.660 4.280 6.800 6.380 ;
        RECT 7.580 4.280 7.720 6.380 ;
        RECT 8.800 5.950 8.940 8.050 ;
        RECT 9.710 5.950 9.850 8.050 ;
        RECT 11.070 7.960 11.580 8.270 ;
        RECT 11.070 6.690 11.210 7.960 ;
        RECT 12.410 6.690 12.550 9.200 ;
        RECT 13.330 6.690 13.470 9.200 ;
        RECT 14.550 8.360 14.690 10.870 ;
        RECT 15.460 8.360 15.600 10.870 ;
        RECT 16.820 10.780 17.330 11.090 ;
        RECT 16.820 9.510 16.960 10.780 ;
        RECT 18.160 9.510 18.300 11.610 ;
        RECT 19.080 9.510 19.220 11.610 ;
        RECT 20.300 11.180 20.440 13.280 ;
        RECT 21.210 11.180 21.350 13.280 ;
        RECT 22.570 13.190 23.080 13.500 ;
        RECT 22.570 11.920 22.710 13.190 ;
        RECT 23.910 11.920 24.050 14.020 ;
        RECT 24.830 11.920 24.970 14.020 ;
        RECT 26.050 13.590 26.190 15.690 ;
        RECT 26.960 13.590 27.100 15.690 ;
        RECT 28.320 15.600 28.830 15.910 ;
        RECT 28.320 14.330 28.460 15.600 ;
        RECT 29.660 14.330 29.800 16.430 ;
        RECT 30.580 14.330 30.720 16.430 ;
        RECT 31.800 16.000 31.940 18.100 ;
        RECT 32.710 16.000 32.850 18.100 ;
        RECT 34.070 18.010 34.580 18.320 ;
        RECT 34.070 16.740 34.210 18.010 ;
        RECT 35.410 16.740 35.550 18.840 ;
        RECT 36.330 16.740 36.470 18.840 ;
        RECT 37.550 18.410 37.690 20.510 ;
        RECT 38.460 18.410 38.600 20.510 ;
        RECT 39.820 20.420 40.330 20.730 ;
        RECT 39.820 19.150 39.960 20.420 ;
        RECT 41.160 19.150 41.300 21.250 ;
        RECT 42.080 19.150 42.220 21.250 ;
        RECT 43.300 20.820 43.440 22.920 ;
        RECT 44.210 20.820 44.350 22.920 ;
        RECT 45.570 22.830 46.080 23.140 ;
        RECT 45.570 21.560 45.710 22.830 ;
        RECT 46.910 21.560 47.050 23.660 ;
        RECT 47.830 21.560 47.970 23.660 ;
        RECT 49.050 23.230 49.190 25.330 ;
        RECT 49.960 23.230 50.100 25.330 ;
        RECT 51.320 25.240 51.830 25.550 ;
        RECT 51.320 23.970 51.460 25.240 ;
        RECT 52.660 23.970 52.800 26.070 ;
        RECT 53.580 23.970 53.720 26.070 ;
        RECT 54.800 25.640 54.940 27.740 ;
        RECT 55.710 25.640 55.850 27.740 ;
        RECT 57.070 27.650 57.580 27.960 ;
        RECT 57.070 26.380 57.210 27.650 ;
        RECT 58.410 26.380 58.550 28.880 ;
        RECT 59.330 26.380 59.470 28.880 ;
        RECT 60.550 28.050 60.690 30.550 ;
        RECT 61.460 28.050 61.600 30.550 ;
        RECT 62.820 30.460 63.330 30.770 ;
        RECT 62.820 29.190 62.960 30.460 ;
        RECT 64.160 29.190 64.300 31.290 ;
        RECT 65.080 29.190 65.220 31.290 ;
        RECT 66.300 30.860 66.440 32.960 ;
        RECT 67.210 30.860 67.350 32.960 ;
        RECT 68.570 32.870 69.080 33.180 ;
        RECT 68.570 31.600 68.710 32.870 ;
        RECT 69.910 31.600 70.050 33.700 ;
        RECT 70.830 31.600 70.970 33.700 ;
        RECT 72.050 33.270 72.190 35.370 ;
        RECT 72.960 33.270 73.100 35.370 ;
        RECT 74.320 35.280 74.830 35.590 ;
        RECT 74.320 34.010 74.460 35.280 ;
        RECT 75.660 34.010 75.800 36.110 ;
        RECT 76.580 34.010 76.720 36.110 ;
        RECT 77.800 35.680 77.940 37.780 ;
        RECT 78.710 35.680 78.850 37.780 ;
        RECT 80.070 37.690 80.580 38.000 ;
        RECT 80.070 36.420 80.210 37.690 ;
        RECT 81.410 36.420 81.550 38.520 ;
        RECT 82.330 36.420 82.470 38.520 ;
        RECT 83.550 38.090 83.690 40.190 ;
        RECT 84.460 38.090 84.600 40.190 ;
        RECT 85.820 40.100 86.330 40.410 ;
        RECT 85.820 38.830 85.960 40.100 ;
        RECT 87.160 38.830 87.300 40.930 ;
        RECT 88.080 38.830 88.220 40.930 ;
        RECT 89.300 40.500 89.440 42.600 ;
        RECT 90.210 40.500 90.350 42.600 ;
        RECT 91.570 42.510 92.080 42.820 ;
        RECT 91.570 41.240 91.710 42.510 ;
        RECT 92.910 41.240 93.050 43.900 ;
        RECT 93.830 41.240 93.970 43.900 ;
        RECT 91.180 40.930 91.710 41.240 ;
        RECT 92.820 40.930 93.140 41.240 ;
        RECT 93.730 40.930 94.050 41.240 ;
        RECT 89.210 40.190 89.530 40.500 ;
        RECT 90.120 40.190 90.440 40.500 ;
        RECT 91.570 40.410 91.710 40.930 ;
        RECT 85.430 38.520 85.960 38.830 ;
        RECT 87.070 38.520 87.390 38.830 ;
        RECT 87.980 38.520 88.300 38.830 ;
        RECT 83.460 37.780 83.780 38.090 ;
        RECT 84.370 37.780 84.690 38.090 ;
        RECT 85.820 38.000 85.960 38.520 ;
        RECT 79.680 36.110 80.210 36.420 ;
        RECT 81.320 36.110 81.640 36.420 ;
        RECT 82.230 36.110 82.550 36.420 ;
        RECT 77.710 35.370 78.030 35.680 ;
        RECT 78.620 35.370 78.940 35.680 ;
        RECT 80.070 35.590 80.210 36.110 ;
        RECT 73.930 33.700 74.460 34.010 ;
        RECT 75.570 33.700 75.890 34.010 ;
        RECT 76.480 33.700 76.800 34.010 ;
        RECT 71.960 32.960 72.280 33.270 ;
        RECT 72.870 32.960 73.190 33.270 ;
        RECT 74.320 33.180 74.460 33.700 ;
        RECT 68.180 31.290 68.710 31.600 ;
        RECT 69.820 31.290 70.140 31.600 ;
        RECT 70.730 31.290 71.050 31.600 ;
        RECT 66.210 30.550 66.530 30.860 ;
        RECT 67.120 30.550 67.440 30.860 ;
        RECT 68.570 30.770 68.710 31.290 ;
        RECT 62.430 28.880 62.960 29.190 ;
        RECT 64.070 28.880 64.390 29.190 ;
        RECT 64.980 28.880 65.300 29.190 ;
        RECT 60.460 27.740 60.780 28.050 ;
        RECT 61.370 27.740 61.690 28.050 ;
        RECT 62.820 27.960 62.960 28.880 ;
        RECT 56.680 26.070 57.210 26.380 ;
        RECT 58.320 26.070 58.640 26.380 ;
        RECT 59.230 26.070 59.550 26.380 ;
        RECT 54.710 25.330 55.030 25.640 ;
        RECT 55.620 25.330 55.940 25.640 ;
        RECT 57.070 25.550 57.210 26.070 ;
        RECT 50.930 23.660 51.460 23.970 ;
        RECT 52.570 23.660 52.890 23.970 ;
        RECT 53.480 23.660 53.800 23.970 ;
        RECT 48.960 22.920 49.280 23.230 ;
        RECT 49.870 22.920 50.190 23.230 ;
        RECT 51.320 23.140 51.460 23.660 ;
        RECT 45.180 21.250 45.710 21.560 ;
        RECT 46.820 21.250 47.140 21.560 ;
        RECT 47.730 21.250 48.050 21.560 ;
        RECT 43.210 20.510 43.530 20.820 ;
        RECT 44.120 20.510 44.440 20.820 ;
        RECT 45.570 20.730 45.710 21.250 ;
        RECT 39.430 18.840 39.960 19.150 ;
        RECT 41.070 18.840 41.390 19.150 ;
        RECT 41.980 18.840 42.300 19.150 ;
        RECT 37.460 18.100 37.780 18.410 ;
        RECT 38.370 18.100 38.690 18.410 ;
        RECT 39.820 18.320 39.960 18.840 ;
        RECT 33.680 16.430 34.210 16.740 ;
        RECT 35.320 16.430 35.640 16.740 ;
        RECT 36.230 16.430 36.550 16.740 ;
        RECT 31.710 15.690 32.030 16.000 ;
        RECT 32.620 15.690 32.940 16.000 ;
        RECT 34.070 15.910 34.210 16.430 ;
        RECT 27.930 14.020 28.460 14.330 ;
        RECT 29.570 14.020 29.890 14.330 ;
        RECT 30.480 14.020 30.800 14.330 ;
        RECT 25.960 13.280 26.280 13.590 ;
        RECT 26.870 13.280 27.190 13.590 ;
        RECT 28.320 13.500 28.460 14.020 ;
        RECT 22.180 11.610 22.710 11.920 ;
        RECT 23.820 11.610 24.140 11.920 ;
        RECT 24.730 11.610 25.050 11.920 ;
        RECT 20.210 10.870 20.530 11.180 ;
        RECT 21.120 10.870 21.440 11.180 ;
        RECT 22.570 11.090 22.710 11.610 ;
        RECT 16.430 9.200 16.960 9.510 ;
        RECT 18.070 9.200 18.390 9.510 ;
        RECT 18.980 9.200 19.300 9.510 ;
        RECT 14.460 8.050 14.780 8.360 ;
        RECT 15.370 8.050 15.690 8.360 ;
        RECT 16.820 8.270 16.960 9.200 ;
        RECT 10.680 6.380 11.210 6.690 ;
        RECT 12.320 6.380 12.640 6.690 ;
        RECT 13.230 6.380 13.550 6.690 ;
        RECT 8.710 5.640 9.030 5.950 ;
        RECT 9.620 5.640 9.940 5.950 ;
        RECT 11.070 5.860 11.210 6.380 ;
        RECT 4.930 3.970 5.460 4.280 ;
        RECT 6.570 3.970 6.890 4.280 ;
        RECT 7.480 3.970 7.800 4.280 ;
        RECT 2.960 3.230 3.280 3.540 ;
        RECT 3.870 3.230 4.190 3.540 ;
        RECT 5.320 3.450 5.460 3.970 ;
        RECT 1.290 1.190 1.550 1.510 ;
        RECT 1.350 -0.900 1.500 1.190 ;
        RECT 3.050 1.130 3.190 3.230 ;
        RECT 3.960 1.130 4.100 3.230 ;
        RECT 5.320 3.140 5.830 3.450 ;
        RECT 5.320 1.870 5.460 3.140 ;
        RECT 6.660 1.870 6.800 3.970 ;
        RECT 7.580 1.870 7.720 3.970 ;
        RECT 8.800 3.540 8.940 5.640 ;
        RECT 9.710 3.540 9.850 5.640 ;
        RECT 11.070 5.550 11.580 5.860 ;
        RECT 11.070 4.280 11.210 5.550 ;
        RECT 12.410 4.280 12.550 6.380 ;
        RECT 13.330 4.280 13.470 6.380 ;
        RECT 14.550 5.950 14.690 8.050 ;
        RECT 15.460 5.950 15.600 8.050 ;
        RECT 16.820 7.960 17.330 8.270 ;
        RECT 16.820 6.690 16.960 7.960 ;
        RECT 18.160 6.690 18.300 9.200 ;
        RECT 19.080 6.690 19.220 9.200 ;
        RECT 20.300 8.360 20.440 10.870 ;
        RECT 21.210 8.360 21.350 10.870 ;
        RECT 22.570 10.780 23.080 11.090 ;
        RECT 22.570 9.510 22.710 10.780 ;
        RECT 23.910 9.510 24.050 11.610 ;
        RECT 24.830 9.510 24.970 11.610 ;
        RECT 26.050 11.180 26.190 13.280 ;
        RECT 26.960 11.180 27.100 13.280 ;
        RECT 28.320 13.190 28.830 13.500 ;
        RECT 28.320 11.920 28.460 13.190 ;
        RECT 29.660 11.920 29.800 14.020 ;
        RECT 30.580 11.920 30.720 14.020 ;
        RECT 31.800 13.590 31.940 15.690 ;
        RECT 32.710 13.590 32.850 15.690 ;
        RECT 34.070 15.600 34.580 15.910 ;
        RECT 34.070 14.330 34.210 15.600 ;
        RECT 35.410 14.330 35.550 16.430 ;
        RECT 36.330 14.330 36.470 16.430 ;
        RECT 37.550 16.000 37.690 18.100 ;
        RECT 38.460 16.000 38.600 18.100 ;
        RECT 39.820 18.010 40.330 18.320 ;
        RECT 39.820 16.740 39.960 18.010 ;
        RECT 41.160 16.740 41.300 18.840 ;
        RECT 42.080 16.740 42.220 18.840 ;
        RECT 43.300 18.410 43.440 20.510 ;
        RECT 44.210 18.410 44.350 20.510 ;
        RECT 45.570 20.420 46.080 20.730 ;
        RECT 45.570 19.150 45.710 20.420 ;
        RECT 46.910 19.150 47.050 21.250 ;
        RECT 47.830 19.150 47.970 21.250 ;
        RECT 49.050 20.820 49.190 22.920 ;
        RECT 49.960 20.820 50.100 22.920 ;
        RECT 51.320 22.830 51.830 23.140 ;
        RECT 51.320 21.560 51.460 22.830 ;
        RECT 52.660 21.560 52.800 23.660 ;
        RECT 53.580 21.560 53.720 23.660 ;
        RECT 54.800 23.230 54.940 25.330 ;
        RECT 55.710 23.230 55.850 25.330 ;
        RECT 57.070 25.240 57.580 25.550 ;
        RECT 57.070 23.970 57.210 25.240 ;
        RECT 58.410 23.970 58.550 26.070 ;
        RECT 59.330 23.970 59.470 26.070 ;
        RECT 60.550 25.640 60.690 27.740 ;
        RECT 61.460 25.640 61.600 27.740 ;
        RECT 62.820 27.650 63.330 27.960 ;
        RECT 62.820 26.380 62.960 27.650 ;
        RECT 64.160 26.380 64.300 28.880 ;
        RECT 65.080 26.380 65.220 28.880 ;
        RECT 66.300 28.050 66.440 30.550 ;
        RECT 67.210 28.050 67.350 30.550 ;
        RECT 68.570 30.460 69.080 30.770 ;
        RECT 68.570 29.190 68.710 30.460 ;
        RECT 69.910 29.190 70.050 31.290 ;
        RECT 70.830 29.190 70.970 31.290 ;
        RECT 72.050 30.860 72.190 32.960 ;
        RECT 72.960 30.860 73.100 32.960 ;
        RECT 74.320 32.870 74.830 33.180 ;
        RECT 74.320 31.600 74.460 32.870 ;
        RECT 75.660 31.600 75.800 33.700 ;
        RECT 76.580 31.600 76.720 33.700 ;
        RECT 77.800 33.270 77.940 35.370 ;
        RECT 78.710 33.270 78.850 35.370 ;
        RECT 80.070 35.280 80.580 35.590 ;
        RECT 80.070 34.010 80.210 35.280 ;
        RECT 81.410 34.010 81.550 36.110 ;
        RECT 82.330 34.010 82.470 36.110 ;
        RECT 83.550 35.680 83.690 37.780 ;
        RECT 84.460 35.680 84.600 37.780 ;
        RECT 85.820 37.690 86.330 38.000 ;
        RECT 85.820 36.420 85.960 37.690 ;
        RECT 87.160 36.420 87.300 38.520 ;
        RECT 88.080 36.420 88.220 38.520 ;
        RECT 89.300 38.090 89.440 40.190 ;
        RECT 90.210 38.090 90.350 40.190 ;
        RECT 91.570 40.100 92.080 40.410 ;
        RECT 91.570 38.830 91.710 40.100 ;
        RECT 92.910 38.830 93.050 40.930 ;
        RECT 93.830 38.830 93.970 40.930 ;
        RECT 91.180 38.520 91.710 38.830 ;
        RECT 92.820 38.520 93.140 38.830 ;
        RECT 93.730 38.520 94.050 38.830 ;
        RECT 89.210 37.780 89.530 38.090 ;
        RECT 90.120 37.780 90.440 38.090 ;
        RECT 91.570 38.000 91.710 38.520 ;
        RECT 85.430 36.110 85.960 36.420 ;
        RECT 87.070 36.110 87.390 36.420 ;
        RECT 87.980 36.110 88.300 36.420 ;
        RECT 83.460 35.370 83.780 35.680 ;
        RECT 84.370 35.370 84.690 35.680 ;
        RECT 85.820 35.590 85.960 36.110 ;
        RECT 79.680 33.700 80.210 34.010 ;
        RECT 81.320 33.700 81.640 34.010 ;
        RECT 82.230 33.700 82.550 34.010 ;
        RECT 77.710 32.960 78.030 33.270 ;
        RECT 78.620 32.960 78.940 33.270 ;
        RECT 80.070 33.180 80.210 33.700 ;
        RECT 73.930 31.290 74.460 31.600 ;
        RECT 75.570 31.290 75.890 31.600 ;
        RECT 76.480 31.290 76.800 31.600 ;
        RECT 71.960 30.550 72.280 30.860 ;
        RECT 72.870 30.550 73.190 30.860 ;
        RECT 74.320 30.770 74.460 31.290 ;
        RECT 68.180 28.880 68.710 29.190 ;
        RECT 69.820 28.880 70.140 29.190 ;
        RECT 70.730 28.880 71.050 29.190 ;
        RECT 66.210 27.740 66.530 28.050 ;
        RECT 67.120 27.740 67.440 28.050 ;
        RECT 68.570 27.960 68.710 28.880 ;
        RECT 62.430 26.070 62.960 26.380 ;
        RECT 64.070 26.070 64.390 26.380 ;
        RECT 64.980 26.070 65.300 26.380 ;
        RECT 60.460 25.330 60.780 25.640 ;
        RECT 61.370 25.330 61.690 25.640 ;
        RECT 62.820 25.550 62.960 26.070 ;
        RECT 56.680 23.660 57.210 23.970 ;
        RECT 58.320 23.660 58.640 23.970 ;
        RECT 59.230 23.660 59.550 23.970 ;
        RECT 54.710 22.920 55.030 23.230 ;
        RECT 55.620 22.920 55.940 23.230 ;
        RECT 57.070 23.140 57.210 23.660 ;
        RECT 50.930 21.250 51.460 21.560 ;
        RECT 52.570 21.250 52.890 21.560 ;
        RECT 53.480 21.250 53.800 21.560 ;
        RECT 48.960 20.510 49.280 20.820 ;
        RECT 49.870 20.510 50.190 20.820 ;
        RECT 51.320 20.730 51.460 21.250 ;
        RECT 45.180 18.840 45.710 19.150 ;
        RECT 46.820 18.840 47.140 19.150 ;
        RECT 47.730 18.840 48.050 19.150 ;
        RECT 43.210 18.100 43.530 18.410 ;
        RECT 44.120 18.100 44.440 18.410 ;
        RECT 45.570 18.320 45.710 18.840 ;
        RECT 39.430 16.430 39.960 16.740 ;
        RECT 41.070 16.430 41.390 16.740 ;
        RECT 41.980 16.430 42.300 16.740 ;
        RECT 37.460 15.690 37.780 16.000 ;
        RECT 38.370 15.690 38.690 16.000 ;
        RECT 39.820 15.910 39.960 16.430 ;
        RECT 33.680 14.020 34.210 14.330 ;
        RECT 35.320 14.020 35.640 14.330 ;
        RECT 36.230 14.020 36.550 14.330 ;
        RECT 31.710 13.280 32.030 13.590 ;
        RECT 32.620 13.280 32.940 13.590 ;
        RECT 34.070 13.500 34.210 14.020 ;
        RECT 27.930 11.610 28.460 11.920 ;
        RECT 29.570 11.610 29.890 11.920 ;
        RECT 30.480 11.610 30.800 11.920 ;
        RECT 25.960 10.870 26.280 11.180 ;
        RECT 26.870 10.870 27.190 11.180 ;
        RECT 28.320 11.090 28.460 11.610 ;
        RECT 22.180 9.200 22.710 9.510 ;
        RECT 23.820 9.200 24.140 9.510 ;
        RECT 24.730 9.200 25.050 9.510 ;
        RECT 20.210 8.050 20.530 8.360 ;
        RECT 21.120 8.050 21.440 8.360 ;
        RECT 22.570 8.270 22.710 9.200 ;
        RECT 16.430 6.380 16.960 6.690 ;
        RECT 18.070 6.380 18.390 6.690 ;
        RECT 18.980 6.380 19.300 6.690 ;
        RECT 14.460 5.640 14.780 5.950 ;
        RECT 15.370 5.640 15.690 5.950 ;
        RECT 16.820 5.860 16.960 6.380 ;
        RECT 10.680 3.970 11.210 4.280 ;
        RECT 12.320 3.970 12.640 4.280 ;
        RECT 13.230 3.970 13.550 4.280 ;
        RECT 8.710 3.230 9.030 3.540 ;
        RECT 9.620 3.230 9.940 3.540 ;
        RECT 11.070 3.450 11.210 3.970 ;
        RECT 4.930 1.560 5.460 1.870 ;
        RECT 6.570 1.560 6.890 1.870 ;
        RECT 7.480 1.560 7.800 1.870 ;
        RECT 2.960 0.820 3.280 1.130 ;
        RECT 3.870 0.820 4.190 1.130 ;
        RECT 5.320 1.040 5.460 1.560 ;
        RECT 1.260 -1.220 1.580 -0.900 ;
        RECT 1.350 -1.750 1.500 -1.220 ;
        RECT 3.050 -1.280 3.190 0.820 ;
        RECT 3.960 -1.280 4.100 0.820 ;
        RECT 5.320 0.730 5.830 1.040 ;
        RECT 5.320 -0.540 5.460 0.730 ;
        RECT 6.660 -0.540 6.800 1.560 ;
        RECT 7.580 -0.540 7.720 1.560 ;
        RECT 8.800 1.130 8.940 3.230 ;
        RECT 9.710 1.130 9.850 3.230 ;
        RECT 11.070 3.140 11.580 3.450 ;
        RECT 11.070 1.870 11.210 3.140 ;
        RECT 12.410 1.870 12.550 3.970 ;
        RECT 13.330 1.870 13.470 3.970 ;
        RECT 14.550 3.540 14.690 5.640 ;
        RECT 15.460 3.540 15.600 5.640 ;
        RECT 16.820 5.550 17.330 5.860 ;
        RECT 16.820 4.280 16.960 5.550 ;
        RECT 18.160 4.280 18.300 6.380 ;
        RECT 19.080 4.280 19.220 6.380 ;
        RECT 20.300 5.950 20.440 8.050 ;
        RECT 21.210 5.950 21.350 8.050 ;
        RECT 22.570 7.960 23.080 8.270 ;
        RECT 22.570 6.690 22.710 7.960 ;
        RECT 23.910 6.690 24.050 9.200 ;
        RECT 24.830 6.690 24.970 9.200 ;
        RECT 26.050 8.360 26.190 10.870 ;
        RECT 26.960 8.360 27.100 10.870 ;
        RECT 28.320 10.780 28.830 11.090 ;
        RECT 28.320 9.510 28.460 10.780 ;
        RECT 29.660 9.510 29.800 11.610 ;
        RECT 30.580 9.510 30.720 11.610 ;
        RECT 31.800 11.180 31.940 13.280 ;
        RECT 32.710 11.180 32.850 13.280 ;
        RECT 34.070 13.190 34.580 13.500 ;
        RECT 34.070 11.920 34.210 13.190 ;
        RECT 35.410 11.920 35.550 14.020 ;
        RECT 36.330 11.920 36.470 14.020 ;
        RECT 37.550 13.590 37.690 15.690 ;
        RECT 38.460 13.590 38.600 15.690 ;
        RECT 39.820 15.600 40.330 15.910 ;
        RECT 39.820 14.330 39.960 15.600 ;
        RECT 41.160 14.330 41.300 16.430 ;
        RECT 42.080 14.330 42.220 16.430 ;
        RECT 43.300 16.000 43.440 18.100 ;
        RECT 44.210 16.000 44.350 18.100 ;
        RECT 45.570 18.010 46.080 18.320 ;
        RECT 45.570 16.740 45.710 18.010 ;
        RECT 46.910 16.740 47.050 18.840 ;
        RECT 47.830 16.740 47.970 18.840 ;
        RECT 49.050 18.410 49.190 20.510 ;
        RECT 49.960 18.410 50.100 20.510 ;
        RECT 51.320 20.420 51.830 20.730 ;
        RECT 51.320 19.150 51.460 20.420 ;
        RECT 52.660 19.150 52.800 21.250 ;
        RECT 53.580 19.150 53.720 21.250 ;
        RECT 54.800 20.820 54.940 22.920 ;
        RECT 55.710 20.820 55.850 22.920 ;
        RECT 57.070 22.830 57.580 23.140 ;
        RECT 57.070 21.560 57.210 22.830 ;
        RECT 58.410 21.560 58.550 23.660 ;
        RECT 59.330 21.560 59.470 23.660 ;
        RECT 60.550 23.230 60.690 25.330 ;
        RECT 61.460 23.230 61.600 25.330 ;
        RECT 62.820 25.240 63.330 25.550 ;
        RECT 62.820 23.970 62.960 25.240 ;
        RECT 64.160 23.970 64.300 26.070 ;
        RECT 65.080 23.970 65.220 26.070 ;
        RECT 66.300 25.640 66.440 27.740 ;
        RECT 67.210 25.640 67.350 27.740 ;
        RECT 68.570 27.650 69.080 27.960 ;
        RECT 68.570 26.380 68.710 27.650 ;
        RECT 69.910 26.380 70.050 28.880 ;
        RECT 70.830 26.380 70.970 28.880 ;
        RECT 72.050 28.050 72.190 30.550 ;
        RECT 72.960 28.050 73.100 30.550 ;
        RECT 74.320 30.460 74.830 30.770 ;
        RECT 74.320 29.190 74.460 30.460 ;
        RECT 75.660 29.190 75.800 31.290 ;
        RECT 76.580 29.190 76.720 31.290 ;
        RECT 77.800 30.860 77.940 32.960 ;
        RECT 78.710 30.860 78.850 32.960 ;
        RECT 80.070 32.870 80.580 33.180 ;
        RECT 80.070 31.600 80.210 32.870 ;
        RECT 81.410 31.600 81.550 33.700 ;
        RECT 82.330 31.600 82.470 33.700 ;
        RECT 83.550 33.270 83.690 35.370 ;
        RECT 84.460 33.270 84.600 35.370 ;
        RECT 85.820 35.280 86.330 35.590 ;
        RECT 85.820 34.010 85.960 35.280 ;
        RECT 87.160 34.010 87.300 36.110 ;
        RECT 88.080 34.010 88.220 36.110 ;
        RECT 89.300 35.680 89.440 37.780 ;
        RECT 90.210 35.680 90.350 37.780 ;
        RECT 91.570 37.690 92.080 38.000 ;
        RECT 91.570 36.420 91.710 37.690 ;
        RECT 92.910 36.420 93.050 38.520 ;
        RECT 93.830 36.420 93.970 38.520 ;
        RECT 91.180 36.110 91.710 36.420 ;
        RECT 92.820 36.110 93.140 36.420 ;
        RECT 93.730 36.110 94.050 36.420 ;
        RECT 89.210 35.370 89.530 35.680 ;
        RECT 90.120 35.370 90.440 35.680 ;
        RECT 91.570 35.590 91.710 36.110 ;
        RECT 85.430 33.700 85.960 34.010 ;
        RECT 87.070 33.700 87.390 34.010 ;
        RECT 87.980 33.700 88.300 34.010 ;
        RECT 83.460 32.960 83.780 33.270 ;
        RECT 84.370 32.960 84.690 33.270 ;
        RECT 85.820 33.180 85.960 33.700 ;
        RECT 79.680 31.290 80.210 31.600 ;
        RECT 81.320 31.290 81.640 31.600 ;
        RECT 82.230 31.290 82.550 31.600 ;
        RECT 77.710 30.550 78.030 30.860 ;
        RECT 78.620 30.550 78.940 30.860 ;
        RECT 80.070 30.770 80.210 31.290 ;
        RECT 73.930 28.880 74.460 29.190 ;
        RECT 75.570 28.880 75.890 29.190 ;
        RECT 76.480 28.880 76.800 29.190 ;
        RECT 71.960 27.740 72.280 28.050 ;
        RECT 72.870 27.740 73.190 28.050 ;
        RECT 74.320 27.960 74.460 28.880 ;
        RECT 68.180 26.070 68.710 26.380 ;
        RECT 69.820 26.070 70.140 26.380 ;
        RECT 70.730 26.070 71.050 26.380 ;
        RECT 66.210 25.330 66.530 25.640 ;
        RECT 67.120 25.330 67.440 25.640 ;
        RECT 68.570 25.550 68.710 26.070 ;
        RECT 62.430 23.660 62.960 23.970 ;
        RECT 64.070 23.660 64.390 23.970 ;
        RECT 64.980 23.660 65.300 23.970 ;
        RECT 60.460 22.920 60.780 23.230 ;
        RECT 61.370 22.920 61.690 23.230 ;
        RECT 62.820 23.140 62.960 23.660 ;
        RECT 56.680 21.250 57.210 21.560 ;
        RECT 58.320 21.250 58.640 21.560 ;
        RECT 59.230 21.250 59.550 21.560 ;
        RECT 54.710 20.510 55.030 20.820 ;
        RECT 55.620 20.510 55.940 20.820 ;
        RECT 57.070 20.730 57.210 21.250 ;
        RECT 50.930 18.840 51.460 19.150 ;
        RECT 52.570 18.840 52.890 19.150 ;
        RECT 53.480 18.840 53.800 19.150 ;
        RECT 48.960 18.100 49.280 18.410 ;
        RECT 49.870 18.100 50.190 18.410 ;
        RECT 51.320 18.320 51.460 18.840 ;
        RECT 45.180 16.430 45.710 16.740 ;
        RECT 46.820 16.430 47.140 16.740 ;
        RECT 47.730 16.430 48.050 16.740 ;
        RECT 43.210 15.690 43.530 16.000 ;
        RECT 44.120 15.690 44.440 16.000 ;
        RECT 45.570 15.910 45.710 16.430 ;
        RECT 39.430 14.020 39.960 14.330 ;
        RECT 41.070 14.020 41.390 14.330 ;
        RECT 41.980 14.020 42.300 14.330 ;
        RECT 37.460 13.280 37.780 13.590 ;
        RECT 38.370 13.280 38.690 13.590 ;
        RECT 39.820 13.500 39.960 14.020 ;
        RECT 33.680 11.610 34.210 11.920 ;
        RECT 35.320 11.610 35.640 11.920 ;
        RECT 36.230 11.610 36.550 11.920 ;
        RECT 31.710 10.870 32.030 11.180 ;
        RECT 32.620 10.870 32.940 11.180 ;
        RECT 34.070 11.090 34.210 11.610 ;
        RECT 27.930 9.200 28.460 9.510 ;
        RECT 29.570 9.200 29.890 9.510 ;
        RECT 30.480 9.200 30.800 9.510 ;
        RECT 25.960 8.050 26.280 8.360 ;
        RECT 26.870 8.050 27.190 8.360 ;
        RECT 28.320 8.270 28.460 9.200 ;
        RECT 22.180 6.380 22.710 6.690 ;
        RECT 23.820 6.380 24.140 6.690 ;
        RECT 24.730 6.380 25.050 6.690 ;
        RECT 20.210 5.640 20.530 5.950 ;
        RECT 21.120 5.640 21.440 5.950 ;
        RECT 22.570 5.860 22.710 6.380 ;
        RECT 16.430 3.970 16.960 4.280 ;
        RECT 18.070 3.970 18.390 4.280 ;
        RECT 18.980 3.970 19.300 4.280 ;
        RECT 14.460 3.230 14.780 3.540 ;
        RECT 15.370 3.230 15.690 3.540 ;
        RECT 16.820 3.450 16.960 3.970 ;
        RECT 10.680 1.560 11.210 1.870 ;
        RECT 12.320 1.560 12.640 1.870 ;
        RECT 13.230 1.560 13.550 1.870 ;
        RECT 8.710 0.820 9.030 1.130 ;
        RECT 9.620 0.820 9.940 1.130 ;
        RECT 11.070 1.040 11.210 1.560 ;
        RECT 4.930 -0.850 5.460 -0.540 ;
        RECT 6.570 -0.850 6.890 -0.540 ;
        RECT 7.480 -0.850 7.800 -0.540 ;
        RECT 2.960 -1.590 3.280 -1.280 ;
        RECT 3.870 -1.590 4.190 -1.280 ;
        RECT 5.320 -1.370 5.460 -0.850 ;
        RECT 1.260 -2.070 1.580 -1.750 ;
        RECT 1.350 -2.540 1.500 -2.070 ;
        RECT 1.260 -2.860 1.580 -2.540 ;
        RECT 1.350 -3.340 1.500 -2.860 ;
        RECT 1.260 -3.600 1.580 -3.340 ;
        RECT 1.350 -4.130 1.500 -3.600 ;
        RECT 3.050 -3.690 3.190 -1.590 ;
        RECT 3.960 -3.690 4.100 -1.590 ;
        RECT 5.320 -1.680 5.830 -1.370 ;
        RECT 5.320 -2.950 5.460 -1.680 ;
        RECT 6.660 -2.950 6.800 -0.850 ;
        RECT 7.580 -2.950 7.720 -0.850 ;
        RECT 8.800 -1.280 8.940 0.820 ;
        RECT 9.710 -1.280 9.850 0.820 ;
        RECT 11.070 0.730 11.580 1.040 ;
        RECT 11.070 -0.540 11.210 0.730 ;
        RECT 12.410 -0.540 12.550 1.560 ;
        RECT 13.330 -0.540 13.470 1.560 ;
        RECT 14.550 1.130 14.690 3.230 ;
        RECT 15.460 1.130 15.600 3.230 ;
        RECT 16.820 3.140 17.330 3.450 ;
        RECT 16.820 1.870 16.960 3.140 ;
        RECT 18.160 1.870 18.300 3.970 ;
        RECT 19.080 1.870 19.220 3.970 ;
        RECT 20.300 3.540 20.440 5.640 ;
        RECT 21.210 3.540 21.350 5.640 ;
        RECT 22.570 5.550 23.080 5.860 ;
        RECT 22.570 4.280 22.710 5.550 ;
        RECT 23.910 4.280 24.050 6.380 ;
        RECT 24.830 4.280 24.970 6.380 ;
        RECT 26.050 5.950 26.190 8.050 ;
        RECT 26.960 5.950 27.100 8.050 ;
        RECT 28.320 7.960 28.830 8.270 ;
        RECT 28.320 6.690 28.460 7.960 ;
        RECT 29.660 6.690 29.800 9.200 ;
        RECT 30.580 6.690 30.720 9.200 ;
        RECT 31.800 8.360 31.940 10.870 ;
        RECT 32.710 8.360 32.850 10.870 ;
        RECT 34.070 10.780 34.580 11.090 ;
        RECT 34.070 9.510 34.210 10.780 ;
        RECT 35.410 9.510 35.550 11.610 ;
        RECT 36.330 9.510 36.470 11.610 ;
        RECT 37.550 11.180 37.690 13.280 ;
        RECT 38.460 11.180 38.600 13.280 ;
        RECT 39.820 13.190 40.330 13.500 ;
        RECT 39.820 11.920 39.960 13.190 ;
        RECT 41.160 11.920 41.300 14.020 ;
        RECT 42.080 11.920 42.220 14.020 ;
        RECT 43.300 13.590 43.440 15.690 ;
        RECT 44.210 13.590 44.350 15.690 ;
        RECT 45.570 15.600 46.080 15.910 ;
        RECT 45.570 14.330 45.710 15.600 ;
        RECT 46.910 14.330 47.050 16.430 ;
        RECT 47.830 14.330 47.970 16.430 ;
        RECT 49.050 16.000 49.190 18.100 ;
        RECT 49.960 16.000 50.100 18.100 ;
        RECT 51.320 18.010 51.830 18.320 ;
        RECT 51.320 16.740 51.460 18.010 ;
        RECT 52.660 16.740 52.800 18.840 ;
        RECT 53.580 16.740 53.720 18.840 ;
        RECT 54.800 18.410 54.940 20.510 ;
        RECT 55.710 18.410 55.850 20.510 ;
        RECT 57.070 20.420 57.580 20.730 ;
        RECT 57.070 19.150 57.210 20.420 ;
        RECT 58.410 19.150 58.550 21.250 ;
        RECT 59.330 19.150 59.470 21.250 ;
        RECT 60.550 20.820 60.690 22.920 ;
        RECT 61.460 20.820 61.600 22.920 ;
        RECT 62.820 22.830 63.330 23.140 ;
        RECT 62.820 21.560 62.960 22.830 ;
        RECT 64.160 21.560 64.300 23.660 ;
        RECT 65.080 21.560 65.220 23.660 ;
        RECT 66.300 23.230 66.440 25.330 ;
        RECT 67.210 23.230 67.350 25.330 ;
        RECT 68.570 25.240 69.080 25.550 ;
        RECT 68.570 23.970 68.710 25.240 ;
        RECT 69.910 23.970 70.050 26.070 ;
        RECT 70.830 23.970 70.970 26.070 ;
        RECT 72.050 25.640 72.190 27.740 ;
        RECT 72.960 25.640 73.100 27.740 ;
        RECT 74.320 27.650 74.830 27.960 ;
        RECT 74.320 26.380 74.460 27.650 ;
        RECT 75.660 26.380 75.800 28.880 ;
        RECT 76.580 26.380 76.720 28.880 ;
        RECT 77.800 28.050 77.940 30.550 ;
        RECT 78.710 28.050 78.850 30.550 ;
        RECT 80.070 30.460 80.580 30.770 ;
        RECT 80.070 29.190 80.210 30.460 ;
        RECT 81.410 29.190 81.550 31.290 ;
        RECT 82.330 29.190 82.470 31.290 ;
        RECT 83.550 30.860 83.690 32.960 ;
        RECT 84.460 30.860 84.600 32.960 ;
        RECT 85.820 32.870 86.330 33.180 ;
        RECT 85.820 31.600 85.960 32.870 ;
        RECT 87.160 31.600 87.300 33.700 ;
        RECT 88.080 31.600 88.220 33.700 ;
        RECT 89.300 33.270 89.440 35.370 ;
        RECT 90.210 33.270 90.350 35.370 ;
        RECT 91.570 35.280 92.080 35.590 ;
        RECT 91.570 34.010 91.710 35.280 ;
        RECT 92.910 34.010 93.050 36.110 ;
        RECT 93.830 34.010 93.970 36.110 ;
        RECT 91.180 33.700 91.710 34.010 ;
        RECT 92.820 33.700 93.140 34.010 ;
        RECT 93.730 33.700 94.050 34.010 ;
        RECT 89.210 32.960 89.530 33.270 ;
        RECT 90.120 32.960 90.440 33.270 ;
        RECT 91.570 33.180 91.710 33.700 ;
        RECT 85.430 31.290 85.960 31.600 ;
        RECT 87.070 31.290 87.390 31.600 ;
        RECT 87.980 31.290 88.300 31.600 ;
        RECT 83.460 30.550 83.780 30.860 ;
        RECT 84.370 30.550 84.690 30.860 ;
        RECT 85.820 30.770 85.960 31.290 ;
        RECT 79.680 28.880 80.210 29.190 ;
        RECT 81.320 28.880 81.640 29.190 ;
        RECT 82.230 28.880 82.550 29.190 ;
        RECT 77.710 27.740 78.030 28.050 ;
        RECT 78.620 27.740 78.940 28.050 ;
        RECT 80.070 27.960 80.210 28.880 ;
        RECT 73.930 26.070 74.460 26.380 ;
        RECT 75.570 26.070 75.890 26.380 ;
        RECT 76.480 26.070 76.800 26.380 ;
        RECT 71.960 25.330 72.280 25.640 ;
        RECT 72.870 25.330 73.190 25.640 ;
        RECT 74.320 25.550 74.460 26.070 ;
        RECT 68.180 23.660 68.710 23.970 ;
        RECT 69.820 23.660 70.140 23.970 ;
        RECT 70.730 23.660 71.050 23.970 ;
        RECT 66.210 22.920 66.530 23.230 ;
        RECT 67.120 22.920 67.440 23.230 ;
        RECT 68.570 23.140 68.710 23.660 ;
        RECT 62.430 21.250 62.960 21.560 ;
        RECT 64.070 21.250 64.390 21.560 ;
        RECT 64.980 21.250 65.300 21.560 ;
        RECT 60.460 20.510 60.780 20.820 ;
        RECT 61.370 20.510 61.690 20.820 ;
        RECT 62.820 20.730 62.960 21.250 ;
        RECT 56.680 18.840 57.210 19.150 ;
        RECT 58.320 18.840 58.640 19.150 ;
        RECT 59.230 18.840 59.550 19.150 ;
        RECT 54.710 18.100 55.030 18.410 ;
        RECT 55.620 18.100 55.940 18.410 ;
        RECT 57.070 18.320 57.210 18.840 ;
        RECT 50.930 16.430 51.460 16.740 ;
        RECT 52.570 16.430 52.890 16.740 ;
        RECT 53.480 16.430 53.800 16.740 ;
        RECT 48.960 15.690 49.280 16.000 ;
        RECT 49.870 15.690 50.190 16.000 ;
        RECT 51.320 15.910 51.460 16.430 ;
        RECT 45.180 14.020 45.710 14.330 ;
        RECT 46.820 14.020 47.140 14.330 ;
        RECT 47.730 14.020 48.050 14.330 ;
        RECT 43.210 13.280 43.530 13.590 ;
        RECT 44.120 13.280 44.440 13.590 ;
        RECT 45.570 13.500 45.710 14.020 ;
        RECT 39.430 11.610 39.960 11.920 ;
        RECT 41.070 11.610 41.390 11.920 ;
        RECT 41.980 11.610 42.300 11.920 ;
        RECT 37.460 10.870 37.780 11.180 ;
        RECT 38.370 10.870 38.690 11.180 ;
        RECT 39.820 11.090 39.960 11.610 ;
        RECT 33.680 9.200 34.210 9.510 ;
        RECT 35.320 9.200 35.640 9.510 ;
        RECT 36.230 9.200 36.550 9.510 ;
        RECT 31.710 8.050 32.030 8.360 ;
        RECT 32.620 8.050 32.940 8.360 ;
        RECT 34.070 8.270 34.210 9.200 ;
        RECT 27.930 6.380 28.460 6.690 ;
        RECT 29.570 6.380 29.890 6.690 ;
        RECT 30.480 6.380 30.800 6.690 ;
        RECT 25.960 5.640 26.280 5.950 ;
        RECT 26.870 5.640 27.190 5.950 ;
        RECT 28.320 5.860 28.460 6.380 ;
        RECT 22.180 3.970 22.710 4.280 ;
        RECT 23.820 3.970 24.140 4.280 ;
        RECT 24.730 3.970 25.050 4.280 ;
        RECT 20.210 3.230 20.530 3.540 ;
        RECT 21.120 3.230 21.440 3.540 ;
        RECT 22.570 3.450 22.710 3.970 ;
        RECT 16.430 1.560 16.960 1.870 ;
        RECT 18.070 1.560 18.390 1.870 ;
        RECT 18.980 1.560 19.300 1.870 ;
        RECT 14.460 0.820 14.780 1.130 ;
        RECT 15.370 0.820 15.690 1.130 ;
        RECT 16.820 1.040 16.960 1.560 ;
        RECT 10.680 -0.850 11.210 -0.540 ;
        RECT 12.320 -0.850 12.640 -0.540 ;
        RECT 13.230 -0.850 13.550 -0.540 ;
        RECT 8.710 -1.590 9.030 -1.280 ;
        RECT 9.620 -1.590 9.940 -1.280 ;
        RECT 11.070 -1.370 11.210 -0.850 ;
        RECT 4.930 -3.260 5.460 -2.950 ;
        RECT 6.570 -3.260 6.890 -2.950 ;
        RECT 7.480 -3.260 7.800 -2.950 ;
        RECT 2.960 -4.000 3.280 -3.690 ;
        RECT 3.870 -4.000 4.190 -3.690 ;
        RECT 5.320 -3.780 5.460 -3.260 ;
        RECT 1.260 -4.450 1.580 -4.130 ;
        RECT 1.350 -4.920 1.500 -4.450 ;
        RECT 1.270 -5.240 1.590 -4.920 ;
        RECT 1.350 -5.720 1.500 -5.240 ;
        RECT 1.290 -6.040 1.550 -5.720 ;
        RECT 1.350 -7.150 1.500 -6.040 ;
        RECT 3.050 -6.690 3.190 -4.000 ;
        RECT 3.960 -6.690 4.100 -4.000 ;
        RECT 5.320 -4.090 5.830 -3.780 ;
        RECT 5.320 -5.360 5.460 -4.090 ;
        RECT 6.660 -5.360 6.800 -3.260 ;
        RECT 7.580 -5.360 7.720 -3.260 ;
        RECT 8.800 -3.690 8.940 -1.590 ;
        RECT 9.710 -3.690 9.850 -1.590 ;
        RECT 11.070 -1.680 11.580 -1.370 ;
        RECT 11.070 -2.950 11.210 -1.680 ;
        RECT 12.410 -2.950 12.550 -0.850 ;
        RECT 13.330 -2.950 13.470 -0.850 ;
        RECT 14.550 -1.280 14.690 0.820 ;
        RECT 15.460 -1.280 15.600 0.820 ;
        RECT 16.820 0.730 17.330 1.040 ;
        RECT 16.820 -0.540 16.960 0.730 ;
        RECT 18.160 -0.540 18.300 1.560 ;
        RECT 19.080 -0.540 19.220 1.560 ;
        RECT 20.300 1.130 20.440 3.230 ;
        RECT 21.210 1.130 21.350 3.230 ;
        RECT 22.570 3.140 23.080 3.450 ;
        RECT 22.570 1.870 22.710 3.140 ;
        RECT 23.910 1.870 24.050 3.970 ;
        RECT 24.830 1.870 24.970 3.970 ;
        RECT 26.050 3.540 26.190 5.640 ;
        RECT 26.960 3.540 27.100 5.640 ;
        RECT 28.320 5.550 28.830 5.860 ;
        RECT 28.320 4.280 28.460 5.550 ;
        RECT 29.660 4.280 29.800 6.380 ;
        RECT 30.580 4.280 30.720 6.380 ;
        RECT 31.800 5.950 31.940 8.050 ;
        RECT 32.710 5.950 32.850 8.050 ;
        RECT 34.070 7.960 34.580 8.270 ;
        RECT 34.070 6.690 34.210 7.960 ;
        RECT 35.410 6.690 35.550 9.200 ;
        RECT 36.330 6.690 36.470 9.200 ;
        RECT 37.550 8.360 37.690 10.870 ;
        RECT 38.460 8.360 38.600 10.870 ;
        RECT 39.820 10.780 40.330 11.090 ;
        RECT 39.820 9.510 39.960 10.780 ;
        RECT 41.160 9.510 41.300 11.610 ;
        RECT 42.080 9.510 42.220 11.610 ;
        RECT 43.300 11.180 43.440 13.280 ;
        RECT 44.210 11.180 44.350 13.280 ;
        RECT 45.570 13.190 46.080 13.500 ;
        RECT 45.570 11.920 45.710 13.190 ;
        RECT 46.910 11.920 47.050 14.020 ;
        RECT 47.830 11.920 47.970 14.020 ;
        RECT 49.050 13.590 49.190 15.690 ;
        RECT 49.960 13.590 50.100 15.690 ;
        RECT 51.320 15.600 51.830 15.910 ;
        RECT 51.320 14.330 51.460 15.600 ;
        RECT 52.660 14.330 52.800 16.430 ;
        RECT 53.580 14.330 53.720 16.430 ;
        RECT 54.800 16.000 54.940 18.100 ;
        RECT 55.710 16.000 55.850 18.100 ;
        RECT 57.070 18.010 57.580 18.320 ;
        RECT 57.070 16.740 57.210 18.010 ;
        RECT 58.410 16.740 58.550 18.840 ;
        RECT 59.330 16.740 59.470 18.840 ;
        RECT 60.550 18.410 60.690 20.510 ;
        RECT 61.460 18.410 61.600 20.510 ;
        RECT 62.820 20.420 63.330 20.730 ;
        RECT 62.820 19.150 62.960 20.420 ;
        RECT 64.160 19.150 64.300 21.250 ;
        RECT 65.080 19.150 65.220 21.250 ;
        RECT 66.300 20.820 66.440 22.920 ;
        RECT 67.210 20.820 67.350 22.920 ;
        RECT 68.570 22.830 69.080 23.140 ;
        RECT 68.570 21.560 68.710 22.830 ;
        RECT 69.910 21.560 70.050 23.660 ;
        RECT 70.830 21.560 70.970 23.660 ;
        RECT 72.050 23.230 72.190 25.330 ;
        RECT 72.960 23.230 73.100 25.330 ;
        RECT 74.320 25.240 74.830 25.550 ;
        RECT 74.320 23.970 74.460 25.240 ;
        RECT 75.660 23.970 75.800 26.070 ;
        RECT 76.580 23.970 76.720 26.070 ;
        RECT 77.800 25.640 77.940 27.740 ;
        RECT 78.710 25.640 78.850 27.740 ;
        RECT 80.070 27.650 80.580 27.960 ;
        RECT 80.070 26.380 80.210 27.650 ;
        RECT 81.410 26.380 81.550 28.880 ;
        RECT 82.330 26.380 82.470 28.880 ;
        RECT 83.550 28.050 83.690 30.550 ;
        RECT 84.460 28.050 84.600 30.550 ;
        RECT 85.820 30.460 86.330 30.770 ;
        RECT 85.820 29.190 85.960 30.460 ;
        RECT 87.160 29.190 87.300 31.290 ;
        RECT 88.080 29.190 88.220 31.290 ;
        RECT 89.300 30.860 89.440 32.960 ;
        RECT 90.210 30.860 90.350 32.960 ;
        RECT 91.570 32.870 92.080 33.180 ;
        RECT 91.570 31.600 91.710 32.870 ;
        RECT 92.910 31.600 93.050 33.700 ;
        RECT 93.830 31.600 93.970 33.700 ;
        RECT 91.180 31.290 91.710 31.600 ;
        RECT 92.820 31.290 93.140 31.600 ;
        RECT 93.730 31.290 94.050 31.600 ;
        RECT 89.210 30.550 89.530 30.860 ;
        RECT 90.120 30.550 90.440 30.860 ;
        RECT 91.570 30.770 91.710 31.290 ;
        RECT 85.430 28.880 85.960 29.190 ;
        RECT 87.070 28.880 87.390 29.190 ;
        RECT 87.980 28.880 88.300 29.190 ;
        RECT 83.460 27.740 83.780 28.050 ;
        RECT 84.370 27.740 84.690 28.050 ;
        RECT 85.820 27.960 85.960 28.880 ;
        RECT 79.680 26.070 80.210 26.380 ;
        RECT 81.320 26.070 81.640 26.380 ;
        RECT 82.230 26.070 82.550 26.380 ;
        RECT 77.710 25.330 78.030 25.640 ;
        RECT 78.620 25.330 78.940 25.640 ;
        RECT 80.070 25.550 80.210 26.070 ;
        RECT 73.930 23.660 74.460 23.970 ;
        RECT 75.570 23.660 75.890 23.970 ;
        RECT 76.480 23.660 76.800 23.970 ;
        RECT 71.960 22.920 72.280 23.230 ;
        RECT 72.870 22.920 73.190 23.230 ;
        RECT 74.320 23.140 74.460 23.660 ;
        RECT 68.180 21.250 68.710 21.560 ;
        RECT 69.820 21.250 70.140 21.560 ;
        RECT 70.730 21.250 71.050 21.560 ;
        RECT 66.210 20.510 66.530 20.820 ;
        RECT 67.120 20.510 67.440 20.820 ;
        RECT 68.570 20.730 68.710 21.250 ;
        RECT 62.430 18.840 62.960 19.150 ;
        RECT 64.070 18.840 64.390 19.150 ;
        RECT 64.980 18.840 65.300 19.150 ;
        RECT 60.460 18.100 60.780 18.410 ;
        RECT 61.370 18.100 61.690 18.410 ;
        RECT 62.820 18.320 62.960 18.840 ;
        RECT 56.680 16.430 57.210 16.740 ;
        RECT 58.320 16.430 58.640 16.740 ;
        RECT 59.230 16.430 59.550 16.740 ;
        RECT 54.710 15.690 55.030 16.000 ;
        RECT 55.620 15.690 55.940 16.000 ;
        RECT 57.070 15.910 57.210 16.430 ;
        RECT 50.930 14.020 51.460 14.330 ;
        RECT 52.570 14.020 52.890 14.330 ;
        RECT 53.480 14.020 53.800 14.330 ;
        RECT 48.960 13.280 49.280 13.590 ;
        RECT 49.870 13.280 50.190 13.590 ;
        RECT 51.320 13.500 51.460 14.020 ;
        RECT 45.180 11.610 45.710 11.920 ;
        RECT 46.820 11.610 47.140 11.920 ;
        RECT 47.730 11.610 48.050 11.920 ;
        RECT 43.210 10.870 43.530 11.180 ;
        RECT 44.120 10.870 44.440 11.180 ;
        RECT 45.570 11.090 45.710 11.610 ;
        RECT 39.430 9.200 39.960 9.510 ;
        RECT 41.070 9.200 41.390 9.510 ;
        RECT 41.980 9.200 42.300 9.510 ;
        RECT 37.460 8.050 37.780 8.360 ;
        RECT 38.370 8.050 38.690 8.360 ;
        RECT 39.820 8.270 39.960 9.200 ;
        RECT 33.680 6.380 34.210 6.690 ;
        RECT 35.320 6.380 35.640 6.690 ;
        RECT 36.230 6.380 36.550 6.690 ;
        RECT 31.710 5.640 32.030 5.950 ;
        RECT 32.620 5.640 32.940 5.950 ;
        RECT 34.070 5.860 34.210 6.380 ;
        RECT 27.930 3.970 28.460 4.280 ;
        RECT 29.570 3.970 29.890 4.280 ;
        RECT 30.480 3.970 30.800 4.280 ;
        RECT 25.960 3.230 26.280 3.540 ;
        RECT 26.870 3.230 27.190 3.540 ;
        RECT 28.320 3.450 28.460 3.970 ;
        RECT 22.180 1.560 22.710 1.870 ;
        RECT 23.820 1.560 24.140 1.870 ;
        RECT 24.730 1.560 25.050 1.870 ;
        RECT 20.210 0.820 20.530 1.130 ;
        RECT 21.120 0.820 21.440 1.130 ;
        RECT 22.570 1.040 22.710 1.560 ;
        RECT 16.430 -0.850 16.960 -0.540 ;
        RECT 18.070 -0.850 18.390 -0.540 ;
        RECT 18.980 -0.850 19.300 -0.540 ;
        RECT 14.460 -1.590 14.780 -1.280 ;
        RECT 15.370 -1.590 15.690 -1.280 ;
        RECT 16.820 -1.370 16.960 -0.850 ;
        RECT 10.680 -3.260 11.210 -2.950 ;
        RECT 12.320 -3.260 12.640 -2.950 ;
        RECT 13.230 -3.260 13.550 -2.950 ;
        RECT 8.710 -4.000 9.030 -3.690 ;
        RECT 9.620 -4.000 9.940 -3.690 ;
        RECT 11.070 -3.780 11.210 -3.260 ;
        RECT 4.930 -5.670 5.460 -5.360 ;
        RECT 6.570 -5.670 6.890 -5.360 ;
        RECT 7.480 -5.670 7.800 -5.360 ;
        RECT 2.960 -7.000 3.280 -6.690 ;
        RECT 3.870 -7.000 4.190 -6.690 ;
        RECT 5.320 -6.780 5.460 -5.670 ;
        RECT 5.960 -6.420 6.260 -6.020 ;
        RECT 1.260 -7.470 1.580 -7.150 ;
        RECT 1.350 -7.950 1.500 -7.470 ;
        RECT 1.260 -8.270 1.580 -7.950 ;
        RECT 1.350 -8.720 1.500 -8.270 ;
        RECT 1.260 -9.040 1.580 -8.720 ;
        RECT 1.350 -9.520 1.500 -9.040 ;
        RECT 3.050 -9.100 3.190 -7.000 ;
        RECT 3.960 -9.100 4.100 -7.000 ;
        RECT 5.320 -7.090 5.830 -6.780 ;
        RECT 5.320 -8.360 5.460 -7.090 ;
        RECT 4.930 -8.670 5.460 -8.360 ;
        RECT 2.960 -9.410 3.280 -9.100 ;
        RECT 3.870 -9.410 4.190 -9.100 ;
        RECT 5.320 -9.190 5.460 -8.670 ;
        RECT 1.260 -9.840 1.580 -9.520 ;
        RECT 1.350 -10.390 1.500 -9.840 ;
        RECT 1.270 -10.710 1.590 -10.390 ;
        RECT 1.350 -11.130 1.500 -10.710 ;
        RECT 1.290 -11.450 1.550 -11.130 ;
        RECT 1.350 -18.900 1.500 -11.450 ;
        RECT 1.290 -19.220 1.550 -18.900 ;
        RECT -41.800 -20.690 -41.500 -20.290 ;
        RECT -0.400 -20.650 0.000 -20.250 ;
        RECT 1.350 -20.300 1.500 -19.220 ;
        RECT 1.260 -20.620 1.590 -20.300 ;
        RECT -43.140 -30.980 -42.840 -30.580 ;
        RECT -41.720 -43.430 -41.580 -20.690 ;
        RECT 3.050 -22.710 3.190 -9.410 ;
        RECT 3.960 -14.240 4.100 -9.410 ;
        RECT 5.320 -9.500 5.830 -9.190 ;
        RECT 5.320 -10.770 5.460 -9.500 ;
        RECT 4.930 -11.080 5.460 -10.770 ;
        RECT 5.320 -12.590 5.460 -11.080 ;
        RECT 5.230 -12.910 5.550 -12.590 ;
        RECT 3.870 -14.570 4.200 -14.240 ;
        RECT 3.960 -19.890 4.100 -14.570 ;
        RECT 3.960 -20.210 4.380 -19.890 ;
        RECT 5.320 -21.780 5.460 -12.910 ;
        RECT 6.020 -13.830 6.190 -6.420 ;
        RECT 6.660 -8.360 6.800 -5.670 ;
        RECT 7.580 -8.360 7.720 -5.670 ;
        RECT 8.800 -6.690 8.940 -4.000 ;
        RECT 9.710 -6.690 9.850 -4.000 ;
        RECT 11.070 -4.090 11.580 -3.780 ;
        RECT 11.070 -5.360 11.210 -4.090 ;
        RECT 12.410 -5.360 12.550 -3.260 ;
        RECT 13.330 -5.360 13.470 -3.260 ;
        RECT 14.550 -3.690 14.690 -1.590 ;
        RECT 15.460 -3.690 15.600 -1.590 ;
        RECT 16.820 -1.680 17.330 -1.370 ;
        RECT 16.820 -2.950 16.960 -1.680 ;
        RECT 18.160 -2.950 18.300 -0.850 ;
        RECT 19.080 -2.950 19.220 -0.850 ;
        RECT 20.300 -1.280 20.440 0.820 ;
        RECT 21.210 -1.280 21.350 0.820 ;
        RECT 22.570 0.730 23.080 1.040 ;
        RECT 22.570 -0.540 22.710 0.730 ;
        RECT 23.910 -0.540 24.050 1.560 ;
        RECT 24.830 -0.540 24.970 1.560 ;
        RECT 26.050 1.130 26.190 3.230 ;
        RECT 26.960 1.130 27.100 3.230 ;
        RECT 28.320 3.140 28.830 3.450 ;
        RECT 28.320 1.870 28.460 3.140 ;
        RECT 29.660 1.870 29.800 3.970 ;
        RECT 30.580 1.870 30.720 3.970 ;
        RECT 31.800 3.540 31.940 5.640 ;
        RECT 32.710 3.540 32.850 5.640 ;
        RECT 34.070 5.550 34.580 5.860 ;
        RECT 34.070 4.280 34.210 5.550 ;
        RECT 35.410 4.280 35.550 6.380 ;
        RECT 36.330 4.280 36.470 6.380 ;
        RECT 37.550 5.950 37.690 8.050 ;
        RECT 38.460 5.950 38.600 8.050 ;
        RECT 39.820 7.960 40.330 8.270 ;
        RECT 39.820 6.690 39.960 7.960 ;
        RECT 41.160 6.690 41.300 9.200 ;
        RECT 42.080 6.690 42.220 9.200 ;
        RECT 43.300 8.360 43.440 10.870 ;
        RECT 44.210 8.360 44.350 10.870 ;
        RECT 45.570 10.780 46.080 11.090 ;
        RECT 45.570 9.510 45.710 10.780 ;
        RECT 46.910 9.510 47.050 11.610 ;
        RECT 47.830 9.510 47.970 11.610 ;
        RECT 49.050 11.180 49.190 13.280 ;
        RECT 49.960 11.180 50.100 13.280 ;
        RECT 51.320 13.190 51.830 13.500 ;
        RECT 51.320 11.920 51.460 13.190 ;
        RECT 52.660 11.920 52.800 14.020 ;
        RECT 53.580 11.920 53.720 14.020 ;
        RECT 54.800 13.590 54.940 15.690 ;
        RECT 55.710 13.590 55.850 15.690 ;
        RECT 57.070 15.600 57.580 15.910 ;
        RECT 57.070 14.330 57.210 15.600 ;
        RECT 58.410 14.330 58.550 16.430 ;
        RECT 59.330 14.330 59.470 16.430 ;
        RECT 60.550 16.000 60.690 18.100 ;
        RECT 61.460 16.000 61.600 18.100 ;
        RECT 62.820 18.010 63.330 18.320 ;
        RECT 62.820 16.740 62.960 18.010 ;
        RECT 64.160 16.740 64.300 18.840 ;
        RECT 65.080 16.740 65.220 18.840 ;
        RECT 66.300 18.410 66.440 20.510 ;
        RECT 67.210 18.410 67.350 20.510 ;
        RECT 68.570 20.420 69.080 20.730 ;
        RECT 68.570 19.150 68.710 20.420 ;
        RECT 69.910 19.150 70.050 21.250 ;
        RECT 70.830 19.150 70.970 21.250 ;
        RECT 72.050 20.820 72.190 22.920 ;
        RECT 72.960 20.820 73.100 22.920 ;
        RECT 74.320 22.830 74.830 23.140 ;
        RECT 74.320 21.560 74.460 22.830 ;
        RECT 75.660 21.560 75.800 23.660 ;
        RECT 76.580 21.560 76.720 23.660 ;
        RECT 77.800 23.230 77.940 25.330 ;
        RECT 78.710 23.230 78.850 25.330 ;
        RECT 80.070 25.240 80.580 25.550 ;
        RECT 80.070 23.970 80.210 25.240 ;
        RECT 81.410 23.970 81.550 26.070 ;
        RECT 82.330 23.970 82.470 26.070 ;
        RECT 83.550 25.640 83.690 27.740 ;
        RECT 84.460 25.640 84.600 27.740 ;
        RECT 85.820 27.650 86.330 27.960 ;
        RECT 85.820 26.380 85.960 27.650 ;
        RECT 87.160 26.380 87.300 28.880 ;
        RECT 88.080 26.380 88.220 28.880 ;
        RECT 89.300 28.050 89.440 30.550 ;
        RECT 90.210 28.050 90.350 30.550 ;
        RECT 91.570 30.460 92.080 30.770 ;
        RECT 91.570 29.190 91.710 30.460 ;
        RECT 92.910 29.190 93.050 31.290 ;
        RECT 93.830 29.190 93.970 31.290 ;
        RECT 91.180 28.880 91.710 29.190 ;
        RECT 92.820 28.880 93.140 29.190 ;
        RECT 93.730 28.880 94.050 29.190 ;
        RECT 89.210 27.740 89.530 28.050 ;
        RECT 90.120 27.740 90.440 28.050 ;
        RECT 91.570 27.960 91.710 28.880 ;
        RECT 85.430 26.070 85.960 26.380 ;
        RECT 87.070 26.070 87.390 26.380 ;
        RECT 87.980 26.070 88.300 26.380 ;
        RECT 83.460 25.330 83.780 25.640 ;
        RECT 84.370 25.330 84.690 25.640 ;
        RECT 85.820 25.550 85.960 26.070 ;
        RECT 79.680 23.660 80.210 23.970 ;
        RECT 81.320 23.660 81.640 23.970 ;
        RECT 82.230 23.660 82.550 23.970 ;
        RECT 77.710 22.920 78.030 23.230 ;
        RECT 78.620 22.920 78.940 23.230 ;
        RECT 80.070 23.140 80.210 23.660 ;
        RECT 73.930 21.250 74.460 21.560 ;
        RECT 75.570 21.250 75.890 21.560 ;
        RECT 76.480 21.250 76.800 21.560 ;
        RECT 71.960 20.510 72.280 20.820 ;
        RECT 72.870 20.510 73.190 20.820 ;
        RECT 74.320 20.730 74.460 21.250 ;
        RECT 68.180 18.840 68.710 19.150 ;
        RECT 69.820 18.840 70.140 19.150 ;
        RECT 70.730 18.840 71.050 19.150 ;
        RECT 66.210 18.100 66.530 18.410 ;
        RECT 67.120 18.100 67.440 18.410 ;
        RECT 68.570 18.320 68.710 18.840 ;
        RECT 62.430 16.430 62.960 16.740 ;
        RECT 64.070 16.430 64.390 16.740 ;
        RECT 64.980 16.430 65.300 16.740 ;
        RECT 60.460 15.690 60.780 16.000 ;
        RECT 61.370 15.690 61.690 16.000 ;
        RECT 62.820 15.910 62.960 16.430 ;
        RECT 56.680 14.020 57.210 14.330 ;
        RECT 58.320 14.020 58.640 14.330 ;
        RECT 59.230 14.020 59.550 14.330 ;
        RECT 54.710 13.280 55.030 13.590 ;
        RECT 55.620 13.280 55.940 13.590 ;
        RECT 57.070 13.500 57.210 14.020 ;
        RECT 50.930 11.610 51.460 11.920 ;
        RECT 52.570 11.610 52.890 11.920 ;
        RECT 53.480 11.610 53.800 11.920 ;
        RECT 48.960 10.870 49.280 11.180 ;
        RECT 49.870 10.870 50.190 11.180 ;
        RECT 51.320 11.090 51.460 11.610 ;
        RECT 45.180 9.200 45.710 9.510 ;
        RECT 46.820 9.200 47.140 9.510 ;
        RECT 47.730 9.200 48.050 9.510 ;
        RECT 43.210 8.050 43.530 8.360 ;
        RECT 44.120 8.050 44.440 8.360 ;
        RECT 45.570 8.270 45.710 9.200 ;
        RECT 39.430 6.380 39.960 6.690 ;
        RECT 41.070 6.380 41.390 6.690 ;
        RECT 41.980 6.380 42.300 6.690 ;
        RECT 37.460 5.640 37.780 5.950 ;
        RECT 38.370 5.640 38.690 5.950 ;
        RECT 39.820 5.860 39.960 6.380 ;
        RECT 33.680 3.970 34.210 4.280 ;
        RECT 35.320 3.970 35.640 4.280 ;
        RECT 36.230 3.970 36.550 4.280 ;
        RECT 31.710 3.230 32.030 3.540 ;
        RECT 32.620 3.230 32.940 3.540 ;
        RECT 34.070 3.450 34.210 3.970 ;
        RECT 27.930 1.560 28.460 1.870 ;
        RECT 29.570 1.560 29.890 1.870 ;
        RECT 30.480 1.560 30.800 1.870 ;
        RECT 25.960 0.820 26.280 1.130 ;
        RECT 26.870 0.820 27.190 1.130 ;
        RECT 28.320 1.040 28.460 1.560 ;
        RECT 22.180 -0.850 22.710 -0.540 ;
        RECT 23.820 -0.850 24.140 -0.540 ;
        RECT 24.730 -0.850 25.050 -0.540 ;
        RECT 20.210 -1.590 20.530 -1.280 ;
        RECT 21.120 -1.590 21.440 -1.280 ;
        RECT 22.570 -1.370 22.710 -0.850 ;
        RECT 16.430 -3.260 16.960 -2.950 ;
        RECT 18.070 -3.260 18.390 -2.950 ;
        RECT 18.980 -3.260 19.300 -2.950 ;
        RECT 14.460 -4.000 14.780 -3.690 ;
        RECT 15.370 -4.000 15.690 -3.690 ;
        RECT 16.820 -3.780 16.960 -3.260 ;
        RECT 10.680 -5.670 11.210 -5.360 ;
        RECT 12.320 -5.670 12.640 -5.360 ;
        RECT 13.230 -5.670 13.550 -5.360 ;
        RECT 8.710 -7.000 9.030 -6.690 ;
        RECT 9.620 -7.000 9.940 -6.690 ;
        RECT 11.070 -6.780 11.210 -5.670 ;
        RECT 6.570 -8.670 6.890 -8.360 ;
        RECT 7.480 -8.670 7.800 -8.360 ;
        RECT 6.660 -10.770 6.800 -8.670 ;
        RECT 7.580 -10.770 7.720 -8.670 ;
        RECT 8.800 -9.100 8.940 -7.000 ;
        RECT 9.710 -9.100 9.850 -7.000 ;
        RECT 11.070 -7.090 11.580 -6.780 ;
        RECT 11.070 -8.360 11.210 -7.090 ;
        RECT 11.710 -7.690 12.010 -7.290 ;
        RECT 10.680 -8.670 11.210 -8.360 ;
        RECT 8.710 -9.410 9.030 -9.100 ;
        RECT 9.620 -9.410 9.940 -9.100 ;
        RECT 11.070 -9.190 11.210 -8.670 ;
        RECT 6.570 -11.080 6.890 -10.770 ;
        RECT 7.480 -11.080 7.800 -10.770 ;
        RECT 5.940 -14.150 6.260 -13.830 ;
        RECT 6.660 -14.240 6.800 -11.080 ;
        RECT 6.580 -14.570 6.910 -14.240 ;
        RECT 6.660 -19.890 6.800 -14.570 ;
        RECT 6.370 -20.210 6.800 -19.890 ;
        RECT 5.230 -22.100 5.550 -21.780 ;
        RECT 2.960 -23.030 3.280 -22.710 ;
        RECT 5.320 -23.380 5.460 -22.100 ;
        RECT 7.580 -22.710 7.720 -11.080 ;
        RECT 8.800 -22.710 8.940 -9.410 ;
        RECT 9.710 -14.240 9.850 -9.410 ;
        RECT 11.070 -9.500 11.580 -9.190 ;
        RECT 11.070 -10.770 11.210 -9.500 ;
        RECT 10.680 -11.080 11.210 -10.770 ;
        RECT 11.070 -12.590 11.210 -11.080 ;
        RECT 10.980 -12.910 11.300 -12.590 ;
        RECT 9.620 -14.570 9.950 -14.240 ;
        RECT 9.710 -19.890 9.850 -14.570 ;
        RECT 9.710 -20.210 10.130 -19.890 ;
        RECT 11.070 -21.780 11.210 -12.910 ;
        RECT 11.770 -13.840 11.940 -7.690 ;
        RECT 12.410 -8.360 12.550 -5.670 ;
        RECT 13.330 -8.360 13.470 -5.670 ;
        RECT 14.550 -6.690 14.690 -4.000 ;
        RECT 15.460 -6.690 15.600 -4.000 ;
        RECT 16.820 -4.090 17.330 -3.780 ;
        RECT 16.820 -5.360 16.960 -4.090 ;
        RECT 18.160 -5.360 18.300 -3.260 ;
        RECT 19.080 -5.360 19.220 -3.260 ;
        RECT 20.300 -3.690 20.440 -1.590 ;
        RECT 21.210 -3.690 21.350 -1.590 ;
        RECT 22.570 -1.680 23.080 -1.370 ;
        RECT 22.570 -2.950 22.710 -1.680 ;
        RECT 23.910 -2.950 24.050 -0.850 ;
        RECT 24.830 -2.950 24.970 -0.850 ;
        RECT 26.050 -1.280 26.190 0.820 ;
        RECT 26.960 -1.280 27.100 0.820 ;
        RECT 28.320 0.730 28.830 1.040 ;
        RECT 28.320 -0.540 28.460 0.730 ;
        RECT 29.660 -0.540 29.800 1.560 ;
        RECT 30.580 -0.540 30.720 1.560 ;
        RECT 31.800 1.130 31.940 3.230 ;
        RECT 32.710 1.130 32.850 3.230 ;
        RECT 34.070 3.140 34.580 3.450 ;
        RECT 34.070 1.870 34.210 3.140 ;
        RECT 35.410 1.870 35.550 3.970 ;
        RECT 36.330 1.870 36.470 3.970 ;
        RECT 37.550 3.540 37.690 5.640 ;
        RECT 38.460 3.540 38.600 5.640 ;
        RECT 39.820 5.550 40.330 5.860 ;
        RECT 39.820 4.280 39.960 5.550 ;
        RECT 41.160 4.280 41.300 6.380 ;
        RECT 42.080 4.280 42.220 6.380 ;
        RECT 43.300 5.950 43.440 8.050 ;
        RECT 44.210 5.950 44.350 8.050 ;
        RECT 45.570 7.960 46.080 8.270 ;
        RECT 45.570 6.690 45.710 7.960 ;
        RECT 46.910 6.690 47.050 9.200 ;
        RECT 47.830 6.690 47.970 9.200 ;
        RECT 49.050 8.360 49.190 10.870 ;
        RECT 49.960 8.360 50.100 10.870 ;
        RECT 51.320 10.780 51.830 11.090 ;
        RECT 51.320 9.510 51.460 10.780 ;
        RECT 52.660 9.510 52.800 11.610 ;
        RECT 53.580 9.510 53.720 11.610 ;
        RECT 54.800 11.180 54.940 13.280 ;
        RECT 55.710 11.180 55.850 13.280 ;
        RECT 57.070 13.190 57.580 13.500 ;
        RECT 57.070 11.920 57.210 13.190 ;
        RECT 58.410 11.920 58.550 14.020 ;
        RECT 59.330 11.920 59.470 14.020 ;
        RECT 60.550 13.590 60.690 15.690 ;
        RECT 61.460 13.590 61.600 15.690 ;
        RECT 62.820 15.600 63.330 15.910 ;
        RECT 62.820 14.330 62.960 15.600 ;
        RECT 64.160 14.330 64.300 16.430 ;
        RECT 65.080 14.330 65.220 16.430 ;
        RECT 66.300 16.000 66.440 18.100 ;
        RECT 67.210 16.000 67.350 18.100 ;
        RECT 68.570 18.010 69.080 18.320 ;
        RECT 68.570 16.740 68.710 18.010 ;
        RECT 69.910 16.740 70.050 18.840 ;
        RECT 70.830 16.740 70.970 18.840 ;
        RECT 72.050 18.410 72.190 20.510 ;
        RECT 72.960 18.410 73.100 20.510 ;
        RECT 74.320 20.420 74.830 20.730 ;
        RECT 74.320 19.150 74.460 20.420 ;
        RECT 75.660 19.150 75.800 21.250 ;
        RECT 76.580 19.150 76.720 21.250 ;
        RECT 77.800 20.820 77.940 22.920 ;
        RECT 78.710 20.820 78.850 22.920 ;
        RECT 80.070 22.830 80.580 23.140 ;
        RECT 80.070 21.560 80.210 22.830 ;
        RECT 81.410 21.560 81.550 23.660 ;
        RECT 82.330 21.560 82.470 23.660 ;
        RECT 83.550 23.230 83.690 25.330 ;
        RECT 84.460 23.230 84.600 25.330 ;
        RECT 85.820 25.240 86.330 25.550 ;
        RECT 85.820 23.970 85.960 25.240 ;
        RECT 87.160 23.970 87.300 26.070 ;
        RECT 88.080 23.970 88.220 26.070 ;
        RECT 89.300 25.640 89.440 27.740 ;
        RECT 90.210 25.640 90.350 27.740 ;
        RECT 91.570 27.650 92.080 27.960 ;
        RECT 91.570 26.380 91.710 27.650 ;
        RECT 92.910 26.380 93.050 28.880 ;
        RECT 93.830 26.380 93.970 28.880 ;
        RECT 91.180 26.070 91.710 26.380 ;
        RECT 92.820 26.070 93.140 26.380 ;
        RECT 93.730 26.070 94.050 26.380 ;
        RECT 89.210 25.330 89.530 25.640 ;
        RECT 90.120 25.330 90.440 25.640 ;
        RECT 91.570 25.550 91.710 26.070 ;
        RECT 85.430 23.660 85.960 23.970 ;
        RECT 87.070 23.660 87.390 23.970 ;
        RECT 87.980 23.660 88.300 23.970 ;
        RECT 83.460 22.920 83.780 23.230 ;
        RECT 84.370 22.920 84.690 23.230 ;
        RECT 85.820 23.140 85.960 23.660 ;
        RECT 79.680 21.250 80.210 21.560 ;
        RECT 81.320 21.250 81.640 21.560 ;
        RECT 82.230 21.250 82.550 21.560 ;
        RECT 77.710 20.510 78.030 20.820 ;
        RECT 78.620 20.510 78.940 20.820 ;
        RECT 80.070 20.730 80.210 21.250 ;
        RECT 73.930 18.840 74.460 19.150 ;
        RECT 75.570 18.840 75.890 19.150 ;
        RECT 76.480 18.840 76.800 19.150 ;
        RECT 71.960 18.100 72.280 18.410 ;
        RECT 72.870 18.100 73.190 18.410 ;
        RECT 74.320 18.320 74.460 18.840 ;
        RECT 68.180 16.430 68.710 16.740 ;
        RECT 69.820 16.430 70.140 16.740 ;
        RECT 70.730 16.430 71.050 16.740 ;
        RECT 66.210 15.690 66.530 16.000 ;
        RECT 67.120 15.690 67.440 16.000 ;
        RECT 68.570 15.910 68.710 16.430 ;
        RECT 62.430 14.020 62.960 14.330 ;
        RECT 64.070 14.020 64.390 14.330 ;
        RECT 64.980 14.020 65.300 14.330 ;
        RECT 60.460 13.280 60.780 13.590 ;
        RECT 61.370 13.280 61.690 13.590 ;
        RECT 62.820 13.500 62.960 14.020 ;
        RECT 56.680 11.610 57.210 11.920 ;
        RECT 58.320 11.610 58.640 11.920 ;
        RECT 59.230 11.610 59.550 11.920 ;
        RECT 54.710 10.870 55.030 11.180 ;
        RECT 55.620 10.870 55.940 11.180 ;
        RECT 57.070 11.090 57.210 11.610 ;
        RECT 50.930 9.200 51.460 9.510 ;
        RECT 52.570 9.200 52.890 9.510 ;
        RECT 53.480 9.200 53.800 9.510 ;
        RECT 48.960 8.050 49.280 8.360 ;
        RECT 49.870 8.050 50.190 8.360 ;
        RECT 51.320 8.270 51.460 9.200 ;
        RECT 45.180 6.380 45.710 6.690 ;
        RECT 46.820 6.380 47.140 6.690 ;
        RECT 47.730 6.380 48.050 6.690 ;
        RECT 43.210 5.640 43.530 5.950 ;
        RECT 44.120 5.640 44.440 5.950 ;
        RECT 45.570 5.860 45.710 6.380 ;
        RECT 39.430 3.970 39.960 4.280 ;
        RECT 41.070 3.970 41.390 4.280 ;
        RECT 41.980 3.970 42.300 4.280 ;
        RECT 37.460 3.230 37.780 3.540 ;
        RECT 38.370 3.230 38.690 3.540 ;
        RECT 39.820 3.450 39.960 3.970 ;
        RECT 33.680 1.560 34.210 1.870 ;
        RECT 35.320 1.560 35.640 1.870 ;
        RECT 36.230 1.560 36.550 1.870 ;
        RECT 31.710 0.820 32.030 1.130 ;
        RECT 32.620 0.820 32.940 1.130 ;
        RECT 34.070 1.040 34.210 1.560 ;
        RECT 27.930 -0.850 28.460 -0.540 ;
        RECT 29.570 -0.850 29.890 -0.540 ;
        RECT 30.480 -0.850 30.800 -0.540 ;
        RECT 25.960 -1.590 26.280 -1.280 ;
        RECT 26.870 -1.590 27.190 -1.280 ;
        RECT 28.320 -1.370 28.460 -0.850 ;
        RECT 22.180 -3.260 22.710 -2.950 ;
        RECT 23.820 -3.260 24.140 -2.950 ;
        RECT 24.730 -3.260 25.050 -2.950 ;
        RECT 20.210 -4.000 20.530 -3.690 ;
        RECT 21.120 -4.000 21.440 -3.690 ;
        RECT 22.570 -3.780 22.710 -3.260 ;
        RECT 16.430 -5.670 16.960 -5.360 ;
        RECT 18.070 -5.670 18.390 -5.360 ;
        RECT 18.980 -5.670 19.300 -5.360 ;
        RECT 14.460 -7.000 14.780 -6.690 ;
        RECT 15.370 -7.000 15.690 -6.690 ;
        RECT 16.820 -6.780 16.960 -5.670 ;
        RECT 12.320 -8.670 12.640 -8.360 ;
        RECT 13.230 -8.670 13.550 -8.360 ;
        RECT 12.410 -10.770 12.550 -8.670 ;
        RECT 13.330 -10.770 13.470 -8.670 ;
        RECT 14.550 -9.100 14.690 -7.000 ;
        RECT 15.460 -9.100 15.600 -7.000 ;
        RECT 16.820 -7.090 17.330 -6.780 ;
        RECT 16.820 -8.360 16.960 -7.090 ;
        RECT 18.160 -8.360 18.300 -5.670 ;
        RECT 19.080 -8.360 19.220 -5.670 ;
        RECT 20.300 -6.690 20.440 -4.000 ;
        RECT 21.210 -6.690 21.350 -4.000 ;
        RECT 22.570 -4.090 23.080 -3.780 ;
        RECT 22.570 -5.360 22.710 -4.090 ;
        RECT 23.910 -5.360 24.050 -3.260 ;
        RECT 24.830 -5.360 24.970 -3.260 ;
        RECT 26.050 -3.690 26.190 -1.590 ;
        RECT 26.960 -3.690 27.100 -1.590 ;
        RECT 28.320 -1.680 28.830 -1.370 ;
        RECT 28.320 -2.950 28.460 -1.680 ;
        RECT 29.660 -2.950 29.800 -0.850 ;
        RECT 30.580 -2.950 30.720 -0.850 ;
        RECT 31.800 -1.280 31.940 0.820 ;
        RECT 32.710 -1.280 32.850 0.820 ;
        RECT 34.070 0.730 34.580 1.040 ;
        RECT 34.070 -0.540 34.210 0.730 ;
        RECT 35.410 -0.540 35.550 1.560 ;
        RECT 36.330 -0.540 36.470 1.560 ;
        RECT 37.550 1.130 37.690 3.230 ;
        RECT 38.460 1.130 38.600 3.230 ;
        RECT 39.820 3.140 40.330 3.450 ;
        RECT 39.820 1.870 39.960 3.140 ;
        RECT 41.160 1.870 41.300 3.970 ;
        RECT 42.080 1.870 42.220 3.970 ;
        RECT 43.300 3.540 43.440 5.640 ;
        RECT 44.210 3.540 44.350 5.640 ;
        RECT 45.570 5.550 46.080 5.860 ;
        RECT 45.570 4.280 45.710 5.550 ;
        RECT 46.910 4.280 47.050 6.380 ;
        RECT 47.830 4.280 47.970 6.380 ;
        RECT 49.050 5.950 49.190 8.050 ;
        RECT 49.960 5.950 50.100 8.050 ;
        RECT 51.320 7.960 51.830 8.270 ;
        RECT 51.320 6.690 51.460 7.960 ;
        RECT 52.660 6.690 52.800 9.200 ;
        RECT 53.580 6.690 53.720 9.200 ;
        RECT 54.800 8.360 54.940 10.870 ;
        RECT 55.710 8.360 55.850 10.870 ;
        RECT 57.070 10.780 57.580 11.090 ;
        RECT 57.070 9.510 57.210 10.780 ;
        RECT 58.410 9.510 58.550 11.610 ;
        RECT 59.330 9.510 59.470 11.610 ;
        RECT 60.550 11.180 60.690 13.280 ;
        RECT 61.460 11.180 61.600 13.280 ;
        RECT 62.820 13.190 63.330 13.500 ;
        RECT 62.820 11.920 62.960 13.190 ;
        RECT 64.160 11.920 64.300 14.020 ;
        RECT 65.080 11.920 65.220 14.020 ;
        RECT 66.300 13.590 66.440 15.690 ;
        RECT 67.210 13.590 67.350 15.690 ;
        RECT 68.570 15.600 69.080 15.910 ;
        RECT 68.570 14.330 68.710 15.600 ;
        RECT 69.910 14.330 70.050 16.430 ;
        RECT 70.830 14.330 70.970 16.430 ;
        RECT 72.050 16.000 72.190 18.100 ;
        RECT 72.960 16.000 73.100 18.100 ;
        RECT 74.320 18.010 74.830 18.320 ;
        RECT 74.320 16.740 74.460 18.010 ;
        RECT 75.660 16.740 75.800 18.840 ;
        RECT 76.580 16.740 76.720 18.840 ;
        RECT 77.800 18.410 77.940 20.510 ;
        RECT 78.710 18.410 78.850 20.510 ;
        RECT 80.070 20.420 80.580 20.730 ;
        RECT 80.070 19.150 80.210 20.420 ;
        RECT 81.410 19.150 81.550 21.250 ;
        RECT 82.330 19.150 82.470 21.250 ;
        RECT 83.550 20.820 83.690 22.920 ;
        RECT 84.460 20.820 84.600 22.920 ;
        RECT 85.820 22.830 86.330 23.140 ;
        RECT 85.820 21.560 85.960 22.830 ;
        RECT 87.160 21.560 87.300 23.660 ;
        RECT 88.080 21.560 88.220 23.660 ;
        RECT 89.300 23.230 89.440 25.330 ;
        RECT 90.210 23.230 90.350 25.330 ;
        RECT 91.570 25.240 92.080 25.550 ;
        RECT 91.570 23.970 91.710 25.240 ;
        RECT 92.910 23.970 93.050 26.070 ;
        RECT 93.830 23.970 93.970 26.070 ;
        RECT 91.180 23.660 91.710 23.970 ;
        RECT 92.820 23.660 93.140 23.970 ;
        RECT 93.730 23.660 94.050 23.970 ;
        RECT 89.210 22.920 89.530 23.230 ;
        RECT 90.120 22.920 90.440 23.230 ;
        RECT 91.570 23.140 91.710 23.660 ;
        RECT 85.430 21.250 85.960 21.560 ;
        RECT 87.070 21.250 87.390 21.560 ;
        RECT 87.980 21.250 88.300 21.560 ;
        RECT 83.460 20.510 83.780 20.820 ;
        RECT 84.370 20.510 84.690 20.820 ;
        RECT 85.820 20.730 85.960 21.250 ;
        RECT 79.680 18.840 80.210 19.150 ;
        RECT 81.320 18.840 81.640 19.150 ;
        RECT 82.230 18.840 82.550 19.150 ;
        RECT 77.710 18.100 78.030 18.410 ;
        RECT 78.620 18.100 78.940 18.410 ;
        RECT 80.070 18.320 80.210 18.840 ;
        RECT 73.930 16.430 74.460 16.740 ;
        RECT 75.570 16.430 75.890 16.740 ;
        RECT 76.480 16.430 76.800 16.740 ;
        RECT 71.960 15.690 72.280 16.000 ;
        RECT 72.870 15.690 73.190 16.000 ;
        RECT 74.320 15.910 74.460 16.430 ;
        RECT 68.180 14.020 68.710 14.330 ;
        RECT 69.820 14.020 70.140 14.330 ;
        RECT 70.730 14.020 71.050 14.330 ;
        RECT 66.210 13.280 66.530 13.590 ;
        RECT 67.120 13.280 67.440 13.590 ;
        RECT 68.570 13.500 68.710 14.020 ;
        RECT 62.430 11.610 62.960 11.920 ;
        RECT 64.070 11.610 64.390 11.920 ;
        RECT 64.980 11.610 65.300 11.920 ;
        RECT 60.460 10.870 60.780 11.180 ;
        RECT 61.370 10.870 61.690 11.180 ;
        RECT 62.820 11.090 62.960 11.610 ;
        RECT 56.680 9.200 57.210 9.510 ;
        RECT 58.320 9.200 58.640 9.510 ;
        RECT 59.230 9.200 59.550 9.510 ;
        RECT 54.710 8.050 55.030 8.360 ;
        RECT 55.620 8.050 55.940 8.360 ;
        RECT 57.070 8.270 57.210 9.200 ;
        RECT 50.930 6.380 51.460 6.690 ;
        RECT 52.570 6.380 52.890 6.690 ;
        RECT 53.480 6.380 53.800 6.690 ;
        RECT 48.960 5.640 49.280 5.950 ;
        RECT 49.870 5.640 50.190 5.950 ;
        RECT 51.320 5.860 51.460 6.380 ;
        RECT 45.180 3.970 45.710 4.280 ;
        RECT 46.820 3.970 47.140 4.280 ;
        RECT 47.730 3.970 48.050 4.280 ;
        RECT 43.210 3.230 43.530 3.540 ;
        RECT 44.120 3.230 44.440 3.540 ;
        RECT 45.570 3.450 45.710 3.970 ;
        RECT 39.430 1.560 39.960 1.870 ;
        RECT 41.070 1.560 41.390 1.870 ;
        RECT 41.980 1.560 42.300 1.870 ;
        RECT 37.460 0.820 37.780 1.130 ;
        RECT 38.370 0.820 38.690 1.130 ;
        RECT 39.820 1.040 39.960 1.560 ;
        RECT 33.680 -0.850 34.210 -0.540 ;
        RECT 35.320 -0.850 35.640 -0.540 ;
        RECT 36.230 -0.850 36.550 -0.540 ;
        RECT 31.710 -1.590 32.030 -1.280 ;
        RECT 32.620 -1.590 32.940 -1.280 ;
        RECT 34.070 -1.370 34.210 -0.850 ;
        RECT 27.930 -3.260 28.460 -2.950 ;
        RECT 29.570 -3.260 29.890 -2.950 ;
        RECT 30.480 -3.260 30.800 -2.950 ;
        RECT 25.960 -4.000 26.280 -3.690 ;
        RECT 26.870 -4.000 27.190 -3.690 ;
        RECT 28.320 -3.780 28.460 -3.260 ;
        RECT 22.180 -5.670 22.710 -5.360 ;
        RECT 23.820 -5.670 24.140 -5.360 ;
        RECT 24.730 -5.670 25.050 -5.360 ;
        RECT 20.210 -7.000 20.530 -6.690 ;
        RECT 21.120 -7.000 21.440 -6.690 ;
        RECT 22.570 -6.780 22.710 -5.670 ;
        RECT 16.430 -8.670 16.960 -8.360 ;
        RECT 14.460 -9.410 14.780 -9.100 ;
        RECT 15.370 -9.410 15.690 -9.100 ;
        RECT 16.820 -9.190 16.960 -8.670 ;
        RECT 17.510 -9.060 17.810 -8.660 ;
        RECT 18.070 -8.670 18.390 -8.360 ;
        RECT 18.980 -8.670 19.300 -8.360 ;
        RECT 12.320 -11.080 12.640 -10.770 ;
        RECT 13.230 -11.080 13.550 -10.770 ;
        RECT 11.690 -14.160 12.010 -13.840 ;
        RECT 12.410 -14.240 12.550 -11.080 ;
        RECT 12.330 -14.570 12.660 -14.240 ;
        RECT 12.410 -19.890 12.550 -14.570 ;
        RECT 12.120 -20.210 12.550 -19.890 ;
        RECT 10.980 -22.100 11.300 -21.780 ;
        RECT 7.490 -23.030 7.810 -22.710 ;
        RECT 8.710 -23.030 9.030 -22.710 ;
        RECT 5.230 -23.700 5.550 -23.380 ;
        RECT 8.060 -23.550 8.460 -23.150 ;
        RECT 11.070 -23.390 11.210 -22.100 ;
        RECT 13.330 -22.710 13.470 -11.080 ;
        RECT 14.550 -22.710 14.690 -9.410 ;
        RECT 15.460 -14.240 15.600 -9.410 ;
        RECT 16.820 -9.500 17.330 -9.190 ;
        RECT 16.820 -10.770 16.960 -9.500 ;
        RECT 16.430 -11.080 16.960 -10.770 ;
        RECT 16.820 -12.590 16.960 -11.080 ;
        RECT 16.730 -12.910 17.050 -12.590 ;
        RECT 15.370 -14.570 15.700 -14.240 ;
        RECT 15.460 -19.890 15.600 -14.570 ;
        RECT 15.460 -20.210 15.880 -19.890 ;
        RECT 16.820 -21.780 16.960 -12.910 ;
        RECT 17.520 -13.860 17.690 -9.060 ;
        RECT 18.160 -10.770 18.300 -8.670 ;
        RECT 19.080 -10.770 19.220 -8.670 ;
        RECT 20.300 -9.100 20.440 -7.000 ;
        RECT 21.210 -9.100 21.350 -7.000 ;
        RECT 22.570 -7.090 23.080 -6.780 ;
        RECT 22.570 -8.360 22.710 -7.090 ;
        RECT 23.910 -8.360 24.050 -5.670 ;
        RECT 24.830 -8.360 24.970 -5.670 ;
        RECT 26.050 -6.690 26.190 -4.000 ;
        RECT 26.960 -6.690 27.100 -4.000 ;
        RECT 28.320 -4.090 28.830 -3.780 ;
        RECT 28.320 -5.360 28.460 -4.090 ;
        RECT 29.660 -5.360 29.800 -3.260 ;
        RECT 30.580 -5.360 30.720 -3.260 ;
        RECT 31.800 -3.690 31.940 -1.590 ;
        RECT 32.710 -3.690 32.850 -1.590 ;
        RECT 34.070 -1.680 34.580 -1.370 ;
        RECT 34.070 -2.950 34.210 -1.680 ;
        RECT 35.410 -2.950 35.550 -0.850 ;
        RECT 36.330 -2.950 36.470 -0.850 ;
        RECT 37.550 -1.280 37.690 0.820 ;
        RECT 38.460 -1.280 38.600 0.820 ;
        RECT 39.820 0.730 40.330 1.040 ;
        RECT 39.820 -0.540 39.960 0.730 ;
        RECT 41.160 -0.540 41.300 1.560 ;
        RECT 42.080 -0.540 42.220 1.560 ;
        RECT 43.300 1.130 43.440 3.230 ;
        RECT 44.210 1.130 44.350 3.230 ;
        RECT 45.570 3.140 46.080 3.450 ;
        RECT 45.570 1.870 45.710 3.140 ;
        RECT 46.910 1.870 47.050 3.970 ;
        RECT 47.830 1.870 47.970 3.970 ;
        RECT 49.050 3.540 49.190 5.640 ;
        RECT 49.960 3.540 50.100 5.640 ;
        RECT 51.320 5.550 51.830 5.860 ;
        RECT 51.320 4.280 51.460 5.550 ;
        RECT 52.660 4.280 52.800 6.380 ;
        RECT 53.580 4.280 53.720 6.380 ;
        RECT 54.800 5.950 54.940 8.050 ;
        RECT 55.710 5.950 55.850 8.050 ;
        RECT 57.070 7.960 57.580 8.270 ;
        RECT 57.070 6.690 57.210 7.960 ;
        RECT 58.410 6.690 58.550 9.200 ;
        RECT 59.330 6.690 59.470 9.200 ;
        RECT 60.550 8.360 60.690 10.870 ;
        RECT 61.460 8.360 61.600 10.870 ;
        RECT 62.820 10.780 63.330 11.090 ;
        RECT 62.820 9.510 62.960 10.780 ;
        RECT 64.160 9.510 64.300 11.610 ;
        RECT 65.080 9.510 65.220 11.610 ;
        RECT 66.300 11.180 66.440 13.280 ;
        RECT 67.210 11.180 67.350 13.280 ;
        RECT 68.570 13.190 69.080 13.500 ;
        RECT 68.570 11.920 68.710 13.190 ;
        RECT 69.910 11.920 70.050 14.020 ;
        RECT 70.830 11.920 70.970 14.020 ;
        RECT 72.050 13.590 72.190 15.690 ;
        RECT 72.960 13.590 73.100 15.690 ;
        RECT 74.320 15.600 74.830 15.910 ;
        RECT 74.320 14.330 74.460 15.600 ;
        RECT 75.660 14.330 75.800 16.430 ;
        RECT 76.580 14.330 76.720 16.430 ;
        RECT 77.800 16.000 77.940 18.100 ;
        RECT 78.710 16.000 78.850 18.100 ;
        RECT 80.070 18.010 80.580 18.320 ;
        RECT 80.070 16.740 80.210 18.010 ;
        RECT 81.410 16.740 81.550 18.840 ;
        RECT 82.330 16.740 82.470 18.840 ;
        RECT 83.550 18.410 83.690 20.510 ;
        RECT 84.460 18.410 84.600 20.510 ;
        RECT 85.820 20.420 86.330 20.730 ;
        RECT 85.820 19.150 85.960 20.420 ;
        RECT 87.160 19.150 87.300 21.250 ;
        RECT 88.080 19.150 88.220 21.250 ;
        RECT 89.300 20.820 89.440 22.920 ;
        RECT 90.210 20.820 90.350 22.920 ;
        RECT 91.570 22.830 92.080 23.140 ;
        RECT 91.570 21.560 91.710 22.830 ;
        RECT 92.910 21.560 93.050 23.660 ;
        RECT 93.830 21.560 93.970 23.660 ;
        RECT 91.180 21.250 91.710 21.560 ;
        RECT 92.820 21.250 93.140 21.560 ;
        RECT 93.730 21.250 94.050 21.560 ;
        RECT 89.210 20.510 89.530 20.820 ;
        RECT 90.120 20.510 90.440 20.820 ;
        RECT 91.570 20.730 91.710 21.250 ;
        RECT 85.430 18.840 85.960 19.150 ;
        RECT 87.070 18.840 87.390 19.150 ;
        RECT 87.980 18.840 88.300 19.150 ;
        RECT 83.460 18.100 83.780 18.410 ;
        RECT 84.370 18.100 84.690 18.410 ;
        RECT 85.820 18.320 85.960 18.840 ;
        RECT 79.680 16.430 80.210 16.740 ;
        RECT 81.320 16.430 81.640 16.740 ;
        RECT 82.230 16.430 82.550 16.740 ;
        RECT 77.710 15.690 78.030 16.000 ;
        RECT 78.620 15.690 78.940 16.000 ;
        RECT 80.070 15.910 80.210 16.430 ;
        RECT 73.930 14.020 74.460 14.330 ;
        RECT 75.570 14.020 75.890 14.330 ;
        RECT 76.480 14.020 76.800 14.330 ;
        RECT 71.960 13.280 72.280 13.590 ;
        RECT 72.870 13.280 73.190 13.590 ;
        RECT 74.320 13.500 74.460 14.020 ;
        RECT 68.180 11.610 68.710 11.920 ;
        RECT 69.820 11.610 70.140 11.920 ;
        RECT 70.730 11.610 71.050 11.920 ;
        RECT 66.210 10.870 66.530 11.180 ;
        RECT 67.120 10.870 67.440 11.180 ;
        RECT 68.570 11.090 68.710 11.610 ;
        RECT 62.430 9.200 62.960 9.510 ;
        RECT 64.070 9.200 64.390 9.510 ;
        RECT 64.980 9.200 65.300 9.510 ;
        RECT 60.460 8.050 60.780 8.360 ;
        RECT 61.370 8.050 61.690 8.360 ;
        RECT 62.820 8.270 62.960 9.200 ;
        RECT 56.680 6.380 57.210 6.690 ;
        RECT 58.320 6.380 58.640 6.690 ;
        RECT 59.230 6.380 59.550 6.690 ;
        RECT 54.710 5.640 55.030 5.950 ;
        RECT 55.620 5.640 55.940 5.950 ;
        RECT 57.070 5.860 57.210 6.380 ;
        RECT 50.930 3.970 51.460 4.280 ;
        RECT 52.570 3.970 52.890 4.280 ;
        RECT 53.480 3.970 53.800 4.280 ;
        RECT 48.960 3.230 49.280 3.540 ;
        RECT 49.870 3.230 50.190 3.540 ;
        RECT 51.320 3.450 51.460 3.970 ;
        RECT 45.180 1.560 45.710 1.870 ;
        RECT 46.820 1.560 47.140 1.870 ;
        RECT 47.730 1.560 48.050 1.870 ;
        RECT 43.210 0.820 43.530 1.130 ;
        RECT 44.120 0.820 44.440 1.130 ;
        RECT 45.570 1.040 45.710 1.560 ;
        RECT 39.430 -0.850 39.960 -0.540 ;
        RECT 41.070 -0.850 41.390 -0.540 ;
        RECT 41.980 -0.850 42.300 -0.540 ;
        RECT 37.460 -1.590 37.780 -1.280 ;
        RECT 38.370 -1.590 38.690 -1.280 ;
        RECT 39.820 -1.370 39.960 -0.850 ;
        RECT 33.680 -3.260 34.210 -2.950 ;
        RECT 35.320 -3.260 35.640 -2.950 ;
        RECT 36.230 -3.260 36.550 -2.950 ;
        RECT 31.710 -4.000 32.030 -3.690 ;
        RECT 32.620 -4.000 32.940 -3.690 ;
        RECT 34.070 -3.780 34.210 -3.260 ;
        RECT 27.930 -5.670 28.460 -5.360 ;
        RECT 29.570 -5.670 29.890 -5.360 ;
        RECT 30.480 -5.670 30.800 -5.360 ;
        RECT 25.960 -7.000 26.280 -6.690 ;
        RECT 26.870 -7.000 27.190 -6.690 ;
        RECT 28.320 -6.780 28.460 -5.670 ;
        RECT 22.180 -8.670 22.710 -8.360 ;
        RECT 23.820 -8.670 24.140 -8.360 ;
        RECT 24.730 -8.670 25.050 -8.360 ;
        RECT 20.210 -9.410 20.530 -9.100 ;
        RECT 21.120 -9.410 21.440 -9.100 ;
        RECT 22.570 -9.190 22.710 -8.670 ;
        RECT 18.070 -11.080 18.390 -10.770 ;
        RECT 18.980 -11.080 19.300 -10.770 ;
        RECT 17.440 -14.180 17.760 -13.860 ;
        RECT 18.160 -14.240 18.300 -11.080 ;
        RECT 18.080 -14.570 18.410 -14.240 ;
        RECT 18.160 -19.890 18.300 -14.570 ;
        RECT 17.870 -20.210 18.300 -19.890 ;
        RECT 16.730 -22.100 17.050 -21.780 ;
        RECT 13.240 -23.030 13.560 -22.710 ;
        RECT 14.460 -23.030 14.780 -22.710 ;
        RECT 10.980 -23.710 11.300 -23.390 ;
        RECT 16.820 -23.440 16.960 -22.100 ;
        RECT 19.080 -22.710 19.220 -11.080 ;
        RECT 20.300 -22.710 20.440 -9.410 ;
        RECT 21.210 -14.240 21.350 -9.410 ;
        RECT 22.570 -9.500 23.080 -9.190 ;
        RECT 22.570 -10.770 22.710 -9.500 ;
        RECT 23.210 -10.230 23.510 -9.830 ;
        RECT 22.180 -11.080 22.710 -10.770 ;
        RECT 22.570 -12.590 22.710 -11.080 ;
        RECT 22.480 -12.910 22.800 -12.590 ;
        RECT 21.120 -14.570 21.450 -14.240 ;
        RECT 21.210 -19.890 21.350 -14.570 ;
        RECT 21.210 -20.210 21.630 -19.890 ;
        RECT 22.570 -21.780 22.710 -12.910 ;
        RECT 23.270 -13.860 23.440 -10.230 ;
        RECT 23.910 -10.770 24.050 -8.670 ;
        RECT 24.830 -10.770 24.970 -8.670 ;
        RECT 26.050 -9.100 26.190 -7.000 ;
        RECT 26.960 -9.100 27.100 -7.000 ;
        RECT 28.320 -7.090 28.830 -6.780 ;
        RECT 28.320 -8.360 28.460 -7.090 ;
        RECT 29.660 -8.360 29.800 -5.670 ;
        RECT 30.580 -8.360 30.720 -5.670 ;
        RECT 31.800 -6.690 31.940 -4.000 ;
        RECT 32.710 -6.690 32.850 -4.000 ;
        RECT 34.070 -4.090 34.580 -3.780 ;
        RECT 34.070 -5.360 34.210 -4.090 ;
        RECT 35.410 -5.360 35.550 -3.260 ;
        RECT 36.330 -5.360 36.470 -3.260 ;
        RECT 37.550 -3.690 37.690 -1.590 ;
        RECT 38.460 -3.690 38.600 -1.590 ;
        RECT 39.820 -1.680 40.330 -1.370 ;
        RECT 39.820 -2.950 39.960 -1.680 ;
        RECT 41.160 -2.950 41.300 -0.850 ;
        RECT 42.080 -2.950 42.220 -0.850 ;
        RECT 43.300 -1.280 43.440 0.820 ;
        RECT 44.210 -1.280 44.350 0.820 ;
        RECT 45.570 0.730 46.080 1.040 ;
        RECT 45.570 -0.540 45.710 0.730 ;
        RECT 46.910 -0.540 47.050 1.560 ;
        RECT 47.830 -0.540 47.970 1.560 ;
        RECT 49.050 1.130 49.190 3.230 ;
        RECT 49.960 1.130 50.100 3.230 ;
        RECT 51.320 3.140 51.830 3.450 ;
        RECT 51.320 1.870 51.460 3.140 ;
        RECT 52.660 1.870 52.800 3.970 ;
        RECT 53.580 1.870 53.720 3.970 ;
        RECT 54.800 3.540 54.940 5.640 ;
        RECT 55.710 3.540 55.850 5.640 ;
        RECT 57.070 5.550 57.580 5.860 ;
        RECT 57.070 4.280 57.210 5.550 ;
        RECT 58.410 4.280 58.550 6.380 ;
        RECT 59.330 4.280 59.470 6.380 ;
        RECT 60.550 5.950 60.690 8.050 ;
        RECT 61.460 5.950 61.600 8.050 ;
        RECT 62.820 7.960 63.330 8.270 ;
        RECT 62.820 6.690 62.960 7.960 ;
        RECT 64.160 6.690 64.300 9.200 ;
        RECT 65.080 6.690 65.220 9.200 ;
        RECT 66.300 8.360 66.440 10.870 ;
        RECT 67.210 8.360 67.350 10.870 ;
        RECT 68.570 10.780 69.080 11.090 ;
        RECT 68.570 9.510 68.710 10.780 ;
        RECT 69.910 9.510 70.050 11.610 ;
        RECT 70.830 9.510 70.970 11.610 ;
        RECT 72.050 11.180 72.190 13.280 ;
        RECT 72.960 11.180 73.100 13.280 ;
        RECT 74.320 13.190 74.830 13.500 ;
        RECT 74.320 11.920 74.460 13.190 ;
        RECT 75.660 11.920 75.800 14.020 ;
        RECT 76.580 11.920 76.720 14.020 ;
        RECT 77.800 13.590 77.940 15.690 ;
        RECT 78.710 13.590 78.850 15.690 ;
        RECT 80.070 15.600 80.580 15.910 ;
        RECT 80.070 14.330 80.210 15.600 ;
        RECT 81.410 14.330 81.550 16.430 ;
        RECT 82.330 14.330 82.470 16.430 ;
        RECT 83.550 16.000 83.690 18.100 ;
        RECT 84.460 16.000 84.600 18.100 ;
        RECT 85.820 18.010 86.330 18.320 ;
        RECT 85.820 16.740 85.960 18.010 ;
        RECT 87.160 16.740 87.300 18.840 ;
        RECT 88.080 16.740 88.220 18.840 ;
        RECT 89.300 18.410 89.440 20.510 ;
        RECT 90.210 18.410 90.350 20.510 ;
        RECT 91.570 20.420 92.080 20.730 ;
        RECT 91.570 19.150 91.710 20.420 ;
        RECT 92.910 19.150 93.050 21.250 ;
        RECT 93.830 19.150 93.970 21.250 ;
        RECT 91.180 18.840 91.710 19.150 ;
        RECT 92.820 18.840 93.140 19.150 ;
        RECT 93.730 18.840 94.050 19.150 ;
        RECT 89.210 18.100 89.530 18.410 ;
        RECT 90.120 18.100 90.440 18.410 ;
        RECT 91.570 18.320 91.710 18.840 ;
        RECT 85.430 16.430 85.960 16.740 ;
        RECT 87.070 16.430 87.390 16.740 ;
        RECT 87.980 16.430 88.300 16.740 ;
        RECT 83.460 15.690 83.780 16.000 ;
        RECT 84.370 15.690 84.690 16.000 ;
        RECT 85.820 15.910 85.960 16.430 ;
        RECT 79.680 14.020 80.210 14.330 ;
        RECT 81.320 14.020 81.640 14.330 ;
        RECT 82.230 14.020 82.550 14.330 ;
        RECT 77.710 13.280 78.030 13.590 ;
        RECT 78.620 13.280 78.940 13.590 ;
        RECT 80.070 13.500 80.210 14.020 ;
        RECT 73.930 11.610 74.460 11.920 ;
        RECT 75.570 11.610 75.890 11.920 ;
        RECT 76.480 11.610 76.800 11.920 ;
        RECT 71.960 10.870 72.280 11.180 ;
        RECT 72.870 10.870 73.190 11.180 ;
        RECT 74.320 11.090 74.460 11.610 ;
        RECT 68.180 9.200 68.710 9.510 ;
        RECT 69.820 9.200 70.140 9.510 ;
        RECT 70.730 9.200 71.050 9.510 ;
        RECT 66.210 8.050 66.530 8.360 ;
        RECT 67.120 8.050 67.440 8.360 ;
        RECT 68.570 8.270 68.710 9.200 ;
        RECT 62.430 6.380 62.960 6.690 ;
        RECT 64.070 6.380 64.390 6.690 ;
        RECT 64.980 6.380 65.300 6.690 ;
        RECT 60.460 5.640 60.780 5.950 ;
        RECT 61.370 5.640 61.690 5.950 ;
        RECT 62.820 5.860 62.960 6.380 ;
        RECT 56.680 3.970 57.210 4.280 ;
        RECT 58.320 3.970 58.640 4.280 ;
        RECT 59.230 3.970 59.550 4.280 ;
        RECT 54.710 3.230 55.030 3.540 ;
        RECT 55.620 3.230 55.940 3.540 ;
        RECT 57.070 3.450 57.210 3.970 ;
        RECT 50.930 1.560 51.460 1.870 ;
        RECT 52.570 1.560 52.890 1.870 ;
        RECT 53.480 1.560 53.800 1.870 ;
        RECT 48.960 0.820 49.280 1.130 ;
        RECT 49.870 0.820 50.190 1.130 ;
        RECT 51.320 1.040 51.460 1.560 ;
        RECT 45.180 -0.850 45.710 -0.540 ;
        RECT 46.820 -0.850 47.140 -0.540 ;
        RECT 47.730 -0.850 48.050 -0.540 ;
        RECT 43.210 -1.590 43.530 -1.280 ;
        RECT 44.120 -1.590 44.440 -1.280 ;
        RECT 45.570 -1.370 45.710 -0.850 ;
        RECT 39.430 -3.260 39.960 -2.950 ;
        RECT 41.070 -3.260 41.390 -2.950 ;
        RECT 41.980 -3.260 42.300 -2.950 ;
        RECT 37.460 -4.000 37.780 -3.690 ;
        RECT 38.370 -4.000 38.690 -3.690 ;
        RECT 39.820 -3.780 39.960 -3.260 ;
        RECT 33.680 -5.670 34.210 -5.360 ;
        RECT 35.320 -5.670 35.640 -5.360 ;
        RECT 36.230 -5.670 36.550 -5.360 ;
        RECT 31.710 -7.000 32.030 -6.690 ;
        RECT 32.620 -7.000 32.940 -6.690 ;
        RECT 34.070 -6.780 34.210 -5.670 ;
        RECT 27.930 -8.670 28.460 -8.360 ;
        RECT 29.570 -8.670 29.890 -8.360 ;
        RECT 30.480 -8.670 30.800 -8.360 ;
        RECT 25.960 -9.410 26.280 -9.100 ;
        RECT 26.870 -9.410 27.190 -9.100 ;
        RECT 28.320 -9.190 28.460 -8.670 ;
        RECT 23.820 -11.080 24.140 -10.770 ;
        RECT 24.730 -11.080 25.050 -10.770 ;
        RECT 23.190 -14.180 23.510 -13.860 ;
        RECT 23.910 -14.240 24.050 -11.080 ;
        RECT 23.830 -14.570 24.160 -14.240 ;
        RECT 23.910 -19.890 24.050 -14.570 ;
        RECT 23.620 -20.210 24.050 -19.890 ;
        RECT 22.480 -22.100 22.800 -21.780 ;
        RECT 18.990 -23.030 19.310 -22.710 ;
        RECT 20.210 -23.030 20.530 -22.710 ;
        RECT 16.730 -23.760 17.050 -23.440 ;
        RECT 19.550 -23.560 19.950 -23.160 ;
        RECT 22.570 -23.440 22.710 -22.100 ;
        RECT 24.830 -22.710 24.970 -11.080 ;
        RECT 26.050 -22.710 26.190 -9.410 ;
        RECT 26.960 -14.240 27.100 -9.410 ;
        RECT 28.320 -9.500 28.830 -9.190 ;
        RECT 28.320 -10.770 28.460 -9.500 ;
        RECT 29.660 -10.770 29.800 -8.670 ;
        RECT 30.580 -10.770 30.720 -8.670 ;
        RECT 31.800 -9.100 31.940 -7.000 ;
        RECT 32.710 -9.100 32.850 -7.000 ;
        RECT 34.070 -7.090 34.580 -6.780 ;
        RECT 34.070 -8.360 34.210 -7.090 ;
        RECT 35.410 -8.360 35.550 -5.670 ;
        RECT 36.330 -8.360 36.470 -5.670 ;
        RECT 37.550 -6.690 37.690 -4.000 ;
        RECT 38.460 -6.690 38.600 -4.000 ;
        RECT 39.820 -4.090 40.330 -3.780 ;
        RECT 39.820 -5.360 39.960 -4.090 ;
        RECT 41.160 -5.360 41.300 -3.260 ;
        RECT 42.080 -5.360 42.220 -3.260 ;
        RECT 43.300 -3.690 43.440 -1.590 ;
        RECT 44.210 -3.690 44.350 -1.590 ;
        RECT 45.570 -1.680 46.080 -1.370 ;
        RECT 45.570 -2.950 45.710 -1.680 ;
        RECT 46.910 -2.950 47.050 -0.850 ;
        RECT 47.830 -2.950 47.970 -0.850 ;
        RECT 49.050 -1.280 49.190 0.820 ;
        RECT 49.960 -1.280 50.100 0.820 ;
        RECT 51.320 0.730 51.830 1.040 ;
        RECT 51.320 -0.540 51.460 0.730 ;
        RECT 52.660 -0.540 52.800 1.560 ;
        RECT 53.580 -0.540 53.720 1.560 ;
        RECT 54.800 1.130 54.940 3.230 ;
        RECT 55.710 1.130 55.850 3.230 ;
        RECT 57.070 3.140 57.580 3.450 ;
        RECT 57.070 1.870 57.210 3.140 ;
        RECT 58.410 1.870 58.550 3.970 ;
        RECT 59.330 1.870 59.470 3.970 ;
        RECT 60.550 3.540 60.690 5.640 ;
        RECT 61.460 3.540 61.600 5.640 ;
        RECT 62.820 5.550 63.330 5.860 ;
        RECT 62.820 4.280 62.960 5.550 ;
        RECT 64.160 4.280 64.300 6.380 ;
        RECT 65.080 4.280 65.220 6.380 ;
        RECT 66.300 5.950 66.440 8.050 ;
        RECT 67.210 5.950 67.350 8.050 ;
        RECT 68.570 7.960 69.080 8.270 ;
        RECT 68.570 6.690 68.710 7.960 ;
        RECT 69.910 6.690 70.050 9.200 ;
        RECT 70.830 6.690 70.970 9.200 ;
        RECT 72.050 8.360 72.190 10.870 ;
        RECT 72.960 8.360 73.100 10.870 ;
        RECT 74.320 10.780 74.830 11.090 ;
        RECT 74.320 9.510 74.460 10.780 ;
        RECT 75.660 9.510 75.800 11.610 ;
        RECT 76.580 9.510 76.720 11.610 ;
        RECT 77.800 11.180 77.940 13.280 ;
        RECT 78.710 11.180 78.850 13.280 ;
        RECT 80.070 13.190 80.580 13.500 ;
        RECT 80.070 11.920 80.210 13.190 ;
        RECT 81.410 11.920 81.550 14.020 ;
        RECT 82.330 11.920 82.470 14.020 ;
        RECT 83.550 13.590 83.690 15.690 ;
        RECT 84.460 13.590 84.600 15.690 ;
        RECT 85.820 15.600 86.330 15.910 ;
        RECT 85.820 14.330 85.960 15.600 ;
        RECT 87.160 14.330 87.300 16.430 ;
        RECT 88.080 14.330 88.220 16.430 ;
        RECT 89.300 16.000 89.440 18.100 ;
        RECT 90.210 16.000 90.350 18.100 ;
        RECT 91.570 18.010 92.080 18.320 ;
        RECT 91.570 16.740 91.710 18.010 ;
        RECT 92.910 16.740 93.050 18.840 ;
        RECT 93.830 16.740 93.970 18.840 ;
        RECT 91.180 16.430 91.710 16.740 ;
        RECT 92.820 16.430 93.140 16.740 ;
        RECT 93.730 16.430 94.050 16.740 ;
        RECT 89.210 15.690 89.530 16.000 ;
        RECT 90.120 15.690 90.440 16.000 ;
        RECT 91.570 15.910 91.710 16.430 ;
        RECT 85.430 14.020 85.960 14.330 ;
        RECT 87.070 14.020 87.390 14.330 ;
        RECT 87.980 14.020 88.300 14.330 ;
        RECT 83.460 13.280 83.780 13.590 ;
        RECT 84.370 13.280 84.690 13.590 ;
        RECT 85.820 13.500 85.960 14.020 ;
        RECT 79.680 11.610 80.210 11.920 ;
        RECT 81.320 11.610 81.640 11.920 ;
        RECT 82.230 11.610 82.550 11.920 ;
        RECT 77.710 10.870 78.030 11.180 ;
        RECT 78.620 10.870 78.940 11.180 ;
        RECT 80.070 11.090 80.210 11.610 ;
        RECT 73.930 9.200 74.460 9.510 ;
        RECT 75.570 9.200 75.890 9.510 ;
        RECT 76.480 9.200 76.800 9.510 ;
        RECT 71.960 8.050 72.280 8.360 ;
        RECT 72.870 8.050 73.190 8.360 ;
        RECT 74.320 8.270 74.460 9.200 ;
        RECT 68.180 6.380 68.710 6.690 ;
        RECT 69.820 6.380 70.140 6.690 ;
        RECT 70.730 6.380 71.050 6.690 ;
        RECT 66.210 5.640 66.530 5.950 ;
        RECT 67.120 5.640 67.440 5.950 ;
        RECT 68.570 5.860 68.710 6.380 ;
        RECT 62.430 3.970 62.960 4.280 ;
        RECT 64.070 3.970 64.390 4.280 ;
        RECT 64.980 3.970 65.300 4.280 ;
        RECT 60.460 3.230 60.780 3.540 ;
        RECT 61.370 3.230 61.690 3.540 ;
        RECT 62.820 3.450 62.960 3.970 ;
        RECT 56.680 1.560 57.210 1.870 ;
        RECT 58.320 1.560 58.640 1.870 ;
        RECT 59.230 1.560 59.550 1.870 ;
        RECT 54.710 0.820 55.030 1.130 ;
        RECT 55.620 0.820 55.940 1.130 ;
        RECT 57.070 1.040 57.210 1.560 ;
        RECT 50.930 -0.850 51.460 -0.540 ;
        RECT 52.570 -0.850 52.890 -0.540 ;
        RECT 53.480 -0.850 53.800 -0.540 ;
        RECT 48.960 -1.590 49.280 -1.280 ;
        RECT 49.870 -1.590 50.190 -1.280 ;
        RECT 51.320 -1.370 51.460 -0.850 ;
        RECT 45.180 -3.260 45.710 -2.950 ;
        RECT 46.820 -3.260 47.140 -2.950 ;
        RECT 47.730 -3.260 48.050 -2.950 ;
        RECT 43.210 -4.000 43.530 -3.690 ;
        RECT 44.120 -4.000 44.440 -3.690 ;
        RECT 45.570 -3.780 45.710 -3.260 ;
        RECT 39.430 -5.670 39.960 -5.360 ;
        RECT 41.070 -5.670 41.390 -5.360 ;
        RECT 41.980 -5.670 42.300 -5.360 ;
        RECT 37.460 -7.000 37.780 -6.690 ;
        RECT 38.370 -7.000 38.690 -6.690 ;
        RECT 39.820 -6.780 39.960 -5.670 ;
        RECT 33.680 -8.670 34.210 -8.360 ;
        RECT 35.320 -8.670 35.640 -8.360 ;
        RECT 36.230 -8.670 36.550 -8.360 ;
        RECT 31.710 -9.410 32.030 -9.100 ;
        RECT 32.620 -9.410 32.940 -9.100 ;
        RECT 34.070 -9.190 34.210 -8.670 ;
        RECT 27.930 -11.080 28.460 -10.770 ;
        RECT 29.570 -11.080 29.890 -10.770 ;
        RECT 30.480 -11.080 30.800 -10.770 ;
        RECT 28.320 -12.590 28.460 -11.080 ;
        RECT 28.960 -11.480 29.260 -11.080 ;
        RECT 28.230 -12.910 28.550 -12.590 ;
        RECT 26.870 -14.570 27.200 -14.240 ;
        RECT 26.960 -19.890 27.100 -14.570 ;
        RECT 26.960 -20.210 27.380 -19.890 ;
        RECT 28.320 -21.780 28.460 -12.910 ;
        RECT 29.020 -13.840 29.190 -11.480 ;
        RECT 28.940 -14.160 29.260 -13.840 ;
        RECT 29.660 -14.240 29.800 -11.080 ;
        RECT 29.580 -14.570 29.910 -14.240 ;
        RECT 29.660 -19.890 29.800 -14.570 ;
        RECT 29.370 -20.210 29.800 -19.890 ;
        RECT 28.230 -22.100 28.550 -21.780 ;
        RECT 24.740 -23.030 25.060 -22.710 ;
        RECT 25.960 -23.030 26.280 -22.710 ;
        RECT 28.320 -23.440 28.460 -22.100 ;
        RECT 30.580 -22.710 30.720 -11.080 ;
        RECT 31.800 -22.710 31.940 -9.410 ;
        RECT 32.710 -14.240 32.850 -9.410 ;
        RECT 34.070 -9.500 34.580 -9.190 ;
        RECT 34.070 -10.770 34.210 -9.500 ;
        RECT 35.410 -10.770 35.550 -8.670 ;
        RECT 36.330 -10.770 36.470 -8.670 ;
        RECT 37.550 -9.100 37.690 -7.000 ;
        RECT 38.460 -9.100 38.600 -7.000 ;
        RECT 39.820 -7.090 40.330 -6.780 ;
        RECT 39.820 -8.360 39.960 -7.090 ;
        RECT 41.160 -8.360 41.300 -5.670 ;
        RECT 42.080 -8.360 42.220 -5.670 ;
        RECT 43.300 -6.690 43.440 -4.000 ;
        RECT 44.210 -6.690 44.350 -4.000 ;
        RECT 45.570 -4.090 46.080 -3.780 ;
        RECT 45.570 -5.360 45.710 -4.090 ;
        RECT 46.910 -5.360 47.050 -3.260 ;
        RECT 47.830 -5.360 47.970 -3.260 ;
        RECT 49.050 -3.690 49.190 -1.590 ;
        RECT 49.960 -3.690 50.100 -1.590 ;
        RECT 51.320 -1.680 51.830 -1.370 ;
        RECT 51.320 -2.950 51.460 -1.680 ;
        RECT 52.660 -2.950 52.800 -0.850 ;
        RECT 53.580 -2.950 53.720 -0.850 ;
        RECT 54.800 -1.280 54.940 0.820 ;
        RECT 55.710 -1.280 55.850 0.820 ;
        RECT 57.070 0.730 57.580 1.040 ;
        RECT 57.070 -0.540 57.210 0.730 ;
        RECT 58.410 -0.540 58.550 1.560 ;
        RECT 59.330 -0.540 59.470 1.560 ;
        RECT 60.550 1.130 60.690 3.230 ;
        RECT 61.460 1.130 61.600 3.230 ;
        RECT 62.820 3.140 63.330 3.450 ;
        RECT 62.820 1.870 62.960 3.140 ;
        RECT 64.160 1.870 64.300 3.970 ;
        RECT 65.080 1.870 65.220 3.970 ;
        RECT 66.300 3.540 66.440 5.640 ;
        RECT 67.210 3.540 67.350 5.640 ;
        RECT 68.570 5.550 69.080 5.860 ;
        RECT 68.570 4.280 68.710 5.550 ;
        RECT 69.910 4.280 70.050 6.380 ;
        RECT 70.830 4.280 70.970 6.380 ;
        RECT 72.050 5.950 72.190 8.050 ;
        RECT 72.960 5.950 73.100 8.050 ;
        RECT 74.320 7.960 74.830 8.270 ;
        RECT 74.320 6.690 74.460 7.960 ;
        RECT 75.660 6.690 75.800 9.200 ;
        RECT 76.580 6.690 76.720 9.200 ;
        RECT 77.800 8.360 77.940 10.870 ;
        RECT 78.710 8.360 78.850 10.870 ;
        RECT 80.070 10.780 80.580 11.090 ;
        RECT 80.070 9.510 80.210 10.780 ;
        RECT 81.410 9.510 81.550 11.610 ;
        RECT 82.330 9.510 82.470 11.610 ;
        RECT 83.550 11.180 83.690 13.280 ;
        RECT 84.460 11.180 84.600 13.280 ;
        RECT 85.820 13.190 86.330 13.500 ;
        RECT 85.820 11.920 85.960 13.190 ;
        RECT 87.160 11.920 87.300 14.020 ;
        RECT 88.080 11.920 88.220 14.020 ;
        RECT 89.300 13.590 89.440 15.690 ;
        RECT 90.210 13.590 90.350 15.690 ;
        RECT 91.570 15.600 92.080 15.910 ;
        RECT 91.570 14.330 91.710 15.600 ;
        RECT 92.910 14.330 93.050 16.430 ;
        RECT 93.830 14.330 93.970 16.430 ;
        RECT 91.180 14.020 91.710 14.330 ;
        RECT 92.820 14.020 93.140 14.330 ;
        RECT 93.730 14.020 94.050 14.330 ;
        RECT 89.210 13.280 89.530 13.590 ;
        RECT 90.120 13.280 90.440 13.590 ;
        RECT 91.570 13.500 91.710 14.020 ;
        RECT 85.430 11.610 85.960 11.920 ;
        RECT 87.070 11.610 87.390 11.920 ;
        RECT 87.980 11.610 88.300 11.920 ;
        RECT 83.460 10.870 83.780 11.180 ;
        RECT 84.370 10.870 84.690 11.180 ;
        RECT 85.820 11.090 85.960 11.610 ;
        RECT 79.680 9.200 80.210 9.510 ;
        RECT 81.320 9.200 81.640 9.510 ;
        RECT 82.230 9.200 82.550 9.510 ;
        RECT 77.710 8.050 78.030 8.360 ;
        RECT 78.620 8.050 78.940 8.360 ;
        RECT 80.070 8.270 80.210 9.200 ;
        RECT 73.930 6.380 74.460 6.690 ;
        RECT 75.570 6.380 75.890 6.690 ;
        RECT 76.480 6.380 76.800 6.690 ;
        RECT 71.960 5.640 72.280 5.950 ;
        RECT 72.870 5.640 73.190 5.950 ;
        RECT 74.320 5.860 74.460 6.380 ;
        RECT 68.180 3.970 68.710 4.280 ;
        RECT 69.820 3.970 70.140 4.280 ;
        RECT 70.730 3.970 71.050 4.280 ;
        RECT 66.210 3.230 66.530 3.540 ;
        RECT 67.120 3.230 67.440 3.540 ;
        RECT 68.570 3.450 68.710 3.970 ;
        RECT 62.430 1.560 62.960 1.870 ;
        RECT 64.070 1.560 64.390 1.870 ;
        RECT 64.980 1.560 65.300 1.870 ;
        RECT 60.460 0.820 60.780 1.130 ;
        RECT 61.370 0.820 61.690 1.130 ;
        RECT 62.820 1.040 62.960 1.560 ;
        RECT 56.680 -0.850 57.210 -0.540 ;
        RECT 58.320 -0.850 58.640 -0.540 ;
        RECT 59.230 -0.850 59.550 -0.540 ;
        RECT 54.710 -1.590 55.030 -1.280 ;
        RECT 55.620 -1.590 55.940 -1.280 ;
        RECT 57.070 -1.370 57.210 -0.850 ;
        RECT 50.930 -3.260 51.460 -2.950 ;
        RECT 52.570 -3.260 52.890 -2.950 ;
        RECT 53.480 -3.260 53.800 -2.950 ;
        RECT 48.960 -4.000 49.280 -3.690 ;
        RECT 49.870 -4.000 50.190 -3.690 ;
        RECT 51.320 -3.780 51.460 -3.260 ;
        RECT 45.180 -5.670 45.710 -5.360 ;
        RECT 46.820 -5.670 47.140 -5.360 ;
        RECT 47.730 -5.670 48.050 -5.360 ;
        RECT 43.210 -7.000 43.530 -6.690 ;
        RECT 44.120 -7.000 44.440 -6.690 ;
        RECT 45.570 -6.780 45.710 -5.670 ;
        RECT 39.430 -8.670 39.960 -8.360 ;
        RECT 41.070 -8.670 41.390 -8.360 ;
        RECT 41.980 -8.670 42.300 -8.360 ;
        RECT 37.460 -9.410 37.780 -9.100 ;
        RECT 38.370 -9.410 38.690 -9.100 ;
        RECT 39.820 -9.190 39.960 -8.670 ;
        RECT 33.680 -11.080 34.210 -10.770 ;
        RECT 35.320 -11.080 35.640 -10.770 ;
        RECT 36.230 -11.080 36.550 -10.770 ;
        RECT 34.070 -12.590 34.210 -11.080 ;
        RECT 33.980 -12.910 34.300 -12.590 ;
        RECT 32.620 -14.570 32.950 -14.240 ;
        RECT 32.710 -19.890 32.850 -14.570 ;
        RECT 32.710 -20.210 33.130 -19.890 ;
        RECT 34.070 -21.780 34.210 -12.910 ;
        RECT 34.710 -12.930 35.010 -12.530 ;
        RECT 34.770 -13.810 34.940 -12.930 ;
        RECT 34.690 -14.130 35.010 -13.810 ;
        RECT 35.410 -14.240 35.550 -11.080 ;
        RECT 35.330 -14.570 35.660 -14.240 ;
        RECT 35.410 -19.890 35.550 -14.570 ;
        RECT 35.120 -20.210 35.550 -19.890 ;
        RECT 33.980 -22.100 34.300 -21.780 ;
        RECT 30.490 -23.030 30.810 -22.710 ;
        RECT 31.710 -23.030 32.030 -22.710 ;
        RECT 22.480 -23.760 22.800 -23.440 ;
        RECT 28.230 -23.760 28.550 -23.440 ;
        RECT 30.980 -23.570 31.380 -23.170 ;
        RECT 34.070 -23.440 34.210 -22.100 ;
        RECT 36.330 -22.710 36.470 -11.080 ;
        RECT 37.550 -22.710 37.690 -9.410 ;
        RECT 38.460 -14.240 38.600 -9.410 ;
        RECT 39.820 -9.500 40.330 -9.190 ;
        RECT 39.820 -10.770 39.960 -9.500 ;
        RECT 41.160 -10.770 41.300 -8.670 ;
        RECT 42.080 -10.770 42.220 -8.670 ;
        RECT 43.300 -9.100 43.440 -7.000 ;
        RECT 44.210 -9.100 44.350 -7.000 ;
        RECT 45.570 -7.090 46.080 -6.780 ;
        RECT 45.570 -8.360 45.710 -7.090 ;
        RECT 46.910 -8.360 47.050 -5.670 ;
        RECT 47.830 -8.360 47.970 -5.670 ;
        RECT 49.050 -6.690 49.190 -4.000 ;
        RECT 49.960 -6.690 50.100 -4.000 ;
        RECT 51.320 -4.090 51.830 -3.780 ;
        RECT 51.320 -5.360 51.460 -4.090 ;
        RECT 52.660 -5.360 52.800 -3.260 ;
        RECT 53.580 -5.360 53.720 -3.260 ;
        RECT 54.800 -3.690 54.940 -1.590 ;
        RECT 55.710 -3.690 55.850 -1.590 ;
        RECT 57.070 -1.680 57.580 -1.370 ;
        RECT 57.070 -2.950 57.210 -1.680 ;
        RECT 58.410 -2.950 58.550 -0.850 ;
        RECT 59.330 -2.950 59.470 -0.850 ;
        RECT 60.550 -1.280 60.690 0.820 ;
        RECT 61.460 -1.280 61.600 0.820 ;
        RECT 62.820 0.730 63.330 1.040 ;
        RECT 62.820 -0.540 62.960 0.730 ;
        RECT 64.160 -0.540 64.300 1.560 ;
        RECT 65.080 -0.540 65.220 1.560 ;
        RECT 66.300 1.130 66.440 3.230 ;
        RECT 67.210 1.130 67.350 3.230 ;
        RECT 68.570 3.140 69.080 3.450 ;
        RECT 68.570 1.870 68.710 3.140 ;
        RECT 69.910 1.870 70.050 3.970 ;
        RECT 70.830 1.870 70.970 3.970 ;
        RECT 72.050 3.540 72.190 5.640 ;
        RECT 72.960 3.540 73.100 5.640 ;
        RECT 74.320 5.550 74.830 5.860 ;
        RECT 74.320 4.280 74.460 5.550 ;
        RECT 75.660 4.280 75.800 6.380 ;
        RECT 76.580 4.280 76.720 6.380 ;
        RECT 77.800 5.950 77.940 8.050 ;
        RECT 78.710 5.950 78.850 8.050 ;
        RECT 80.070 7.960 80.580 8.270 ;
        RECT 80.070 6.690 80.210 7.960 ;
        RECT 81.410 6.690 81.550 9.200 ;
        RECT 82.330 6.690 82.470 9.200 ;
        RECT 83.550 8.360 83.690 10.870 ;
        RECT 84.460 8.360 84.600 10.870 ;
        RECT 85.820 10.780 86.330 11.090 ;
        RECT 85.820 9.510 85.960 10.780 ;
        RECT 87.160 9.510 87.300 11.610 ;
        RECT 88.080 9.510 88.220 11.610 ;
        RECT 89.300 11.180 89.440 13.280 ;
        RECT 90.210 11.180 90.350 13.280 ;
        RECT 91.570 13.190 92.080 13.500 ;
        RECT 91.570 11.920 91.710 13.190 ;
        RECT 92.910 11.920 93.050 14.020 ;
        RECT 93.830 11.920 93.970 14.020 ;
        RECT 91.180 11.610 91.710 11.920 ;
        RECT 92.820 11.610 93.140 11.920 ;
        RECT 93.730 11.610 94.050 11.920 ;
        RECT 89.210 10.870 89.530 11.180 ;
        RECT 90.120 10.870 90.440 11.180 ;
        RECT 91.570 11.090 91.710 11.610 ;
        RECT 85.430 9.200 85.960 9.510 ;
        RECT 87.070 9.200 87.390 9.510 ;
        RECT 87.980 9.200 88.300 9.510 ;
        RECT 83.460 8.050 83.780 8.360 ;
        RECT 84.370 8.050 84.690 8.360 ;
        RECT 85.820 8.270 85.960 9.200 ;
        RECT 79.680 6.380 80.210 6.690 ;
        RECT 81.320 6.380 81.640 6.690 ;
        RECT 82.230 6.380 82.550 6.690 ;
        RECT 77.710 5.640 78.030 5.950 ;
        RECT 78.620 5.640 78.940 5.950 ;
        RECT 80.070 5.860 80.210 6.380 ;
        RECT 73.930 3.970 74.460 4.280 ;
        RECT 75.570 3.970 75.890 4.280 ;
        RECT 76.480 3.970 76.800 4.280 ;
        RECT 71.960 3.230 72.280 3.540 ;
        RECT 72.870 3.230 73.190 3.540 ;
        RECT 74.320 3.450 74.460 3.970 ;
        RECT 68.180 1.560 68.710 1.870 ;
        RECT 69.820 1.560 70.140 1.870 ;
        RECT 70.730 1.560 71.050 1.870 ;
        RECT 66.210 0.820 66.530 1.130 ;
        RECT 67.120 0.820 67.440 1.130 ;
        RECT 68.570 1.040 68.710 1.560 ;
        RECT 62.430 -0.850 62.960 -0.540 ;
        RECT 64.070 -0.850 64.390 -0.540 ;
        RECT 64.980 -0.850 65.300 -0.540 ;
        RECT 60.460 -1.590 60.780 -1.280 ;
        RECT 61.370 -1.590 61.690 -1.280 ;
        RECT 62.820 -1.370 62.960 -0.850 ;
        RECT 56.680 -3.260 57.210 -2.950 ;
        RECT 58.320 -3.260 58.640 -2.950 ;
        RECT 59.230 -3.260 59.550 -2.950 ;
        RECT 54.710 -4.000 55.030 -3.690 ;
        RECT 55.620 -4.000 55.940 -3.690 ;
        RECT 57.070 -3.780 57.210 -3.260 ;
        RECT 50.930 -5.670 51.460 -5.360 ;
        RECT 52.570 -5.670 52.890 -5.360 ;
        RECT 53.480 -5.670 53.800 -5.360 ;
        RECT 48.960 -7.000 49.280 -6.690 ;
        RECT 49.870 -7.000 50.190 -6.690 ;
        RECT 51.320 -6.780 51.460 -5.670 ;
        RECT 45.180 -8.670 45.710 -8.360 ;
        RECT 46.820 -8.670 47.140 -8.360 ;
        RECT 47.730 -8.670 48.050 -8.360 ;
        RECT 43.210 -9.410 43.530 -9.100 ;
        RECT 44.120 -9.410 44.440 -9.100 ;
        RECT 45.570 -9.190 45.710 -8.670 ;
        RECT 39.430 -11.080 39.960 -10.770 ;
        RECT 41.070 -11.080 41.390 -10.770 ;
        RECT 41.980 -11.080 42.300 -10.770 ;
        RECT 39.820 -12.590 39.960 -11.080 ;
        RECT 39.730 -12.910 40.050 -12.590 ;
        RECT 38.370 -14.570 38.700 -14.240 ;
        RECT 38.460 -19.890 38.600 -14.570 ;
        RECT 38.460 -20.210 38.880 -19.890 ;
        RECT 39.820 -21.780 39.960 -12.910 ;
        RECT 40.400 -14.150 40.800 -13.750 ;
        RECT 41.160 -14.240 41.300 -11.080 ;
        RECT 41.080 -14.570 41.410 -14.240 ;
        RECT 41.160 -19.890 41.300 -14.570 ;
        RECT 40.870 -20.210 41.300 -19.890 ;
        RECT 39.730 -22.100 40.050 -21.780 ;
        RECT 36.240 -23.030 36.560 -22.710 ;
        RECT 37.460 -23.030 37.780 -22.710 ;
        RECT 39.820 -23.440 39.960 -22.100 ;
        RECT 42.080 -22.710 42.220 -11.080 ;
        RECT 43.300 -22.710 43.440 -9.410 ;
        RECT 44.210 -14.240 44.350 -9.410 ;
        RECT 45.570 -9.500 46.080 -9.190 ;
        RECT 45.570 -10.770 45.710 -9.500 ;
        RECT 46.910 -10.770 47.050 -8.670 ;
        RECT 47.830 -10.770 47.970 -8.670 ;
        RECT 49.050 -9.100 49.190 -7.000 ;
        RECT 49.960 -9.100 50.100 -7.000 ;
        RECT 51.320 -7.090 51.830 -6.780 ;
        RECT 51.320 -8.360 51.460 -7.090 ;
        RECT 52.660 -8.360 52.800 -5.670 ;
        RECT 53.580 -8.360 53.720 -5.670 ;
        RECT 54.800 -6.690 54.940 -4.000 ;
        RECT 55.710 -6.690 55.850 -4.000 ;
        RECT 57.070 -4.090 57.580 -3.780 ;
        RECT 57.070 -5.360 57.210 -4.090 ;
        RECT 58.410 -5.360 58.550 -3.260 ;
        RECT 59.330 -5.360 59.470 -3.260 ;
        RECT 60.550 -3.690 60.690 -1.590 ;
        RECT 61.460 -3.690 61.600 -1.590 ;
        RECT 62.820 -1.680 63.330 -1.370 ;
        RECT 62.820 -2.950 62.960 -1.680 ;
        RECT 64.160 -2.950 64.300 -0.850 ;
        RECT 65.080 -2.950 65.220 -0.850 ;
        RECT 66.300 -1.280 66.440 0.820 ;
        RECT 67.210 -1.280 67.350 0.820 ;
        RECT 68.570 0.730 69.080 1.040 ;
        RECT 68.570 -0.540 68.710 0.730 ;
        RECT 69.910 -0.540 70.050 1.560 ;
        RECT 70.830 -0.540 70.970 1.560 ;
        RECT 72.050 1.130 72.190 3.230 ;
        RECT 72.960 1.130 73.100 3.230 ;
        RECT 74.320 3.140 74.830 3.450 ;
        RECT 74.320 1.870 74.460 3.140 ;
        RECT 75.660 1.870 75.800 3.970 ;
        RECT 76.580 1.870 76.720 3.970 ;
        RECT 77.800 3.540 77.940 5.640 ;
        RECT 78.710 3.540 78.850 5.640 ;
        RECT 80.070 5.550 80.580 5.860 ;
        RECT 80.070 4.280 80.210 5.550 ;
        RECT 81.410 4.280 81.550 6.380 ;
        RECT 82.330 4.280 82.470 6.380 ;
        RECT 83.550 5.950 83.690 8.050 ;
        RECT 84.460 5.950 84.600 8.050 ;
        RECT 85.820 7.960 86.330 8.270 ;
        RECT 85.820 6.690 85.960 7.960 ;
        RECT 87.160 6.690 87.300 9.200 ;
        RECT 88.080 6.690 88.220 9.200 ;
        RECT 89.300 8.360 89.440 10.870 ;
        RECT 90.210 8.360 90.350 10.870 ;
        RECT 91.570 10.780 92.080 11.090 ;
        RECT 91.570 9.510 91.710 10.780 ;
        RECT 92.910 9.510 93.050 11.610 ;
        RECT 93.830 9.510 93.970 11.610 ;
        RECT 91.180 9.200 91.710 9.510 ;
        RECT 92.820 9.200 93.140 9.510 ;
        RECT 93.730 9.200 94.050 9.510 ;
        RECT 89.210 8.050 89.530 8.360 ;
        RECT 90.120 8.050 90.440 8.360 ;
        RECT 91.570 8.270 91.710 9.200 ;
        RECT 85.430 6.380 85.960 6.690 ;
        RECT 87.070 6.380 87.390 6.690 ;
        RECT 87.980 6.380 88.300 6.690 ;
        RECT 83.460 5.640 83.780 5.950 ;
        RECT 84.370 5.640 84.690 5.950 ;
        RECT 85.820 5.860 85.960 6.380 ;
        RECT 79.680 3.970 80.210 4.280 ;
        RECT 81.320 3.970 81.640 4.280 ;
        RECT 82.230 3.970 82.550 4.280 ;
        RECT 77.710 3.230 78.030 3.540 ;
        RECT 78.620 3.230 78.940 3.540 ;
        RECT 80.070 3.450 80.210 3.970 ;
        RECT 73.930 1.560 74.460 1.870 ;
        RECT 75.570 1.560 75.890 1.870 ;
        RECT 76.480 1.560 76.800 1.870 ;
        RECT 71.960 0.820 72.280 1.130 ;
        RECT 72.870 0.820 73.190 1.130 ;
        RECT 74.320 1.040 74.460 1.560 ;
        RECT 68.180 -0.850 68.710 -0.540 ;
        RECT 69.820 -0.850 70.140 -0.540 ;
        RECT 70.730 -0.850 71.050 -0.540 ;
        RECT 66.210 -1.590 66.530 -1.280 ;
        RECT 67.120 -1.590 67.440 -1.280 ;
        RECT 68.570 -1.370 68.710 -0.850 ;
        RECT 62.430 -3.260 62.960 -2.950 ;
        RECT 64.070 -3.260 64.390 -2.950 ;
        RECT 64.980 -3.260 65.300 -2.950 ;
        RECT 60.460 -4.000 60.780 -3.690 ;
        RECT 61.370 -4.000 61.690 -3.690 ;
        RECT 62.820 -3.780 62.960 -3.260 ;
        RECT 56.680 -5.670 57.210 -5.360 ;
        RECT 58.320 -5.670 58.640 -5.360 ;
        RECT 59.230 -5.670 59.550 -5.360 ;
        RECT 54.710 -7.000 55.030 -6.690 ;
        RECT 55.620 -7.000 55.940 -6.690 ;
        RECT 57.070 -6.780 57.210 -5.670 ;
        RECT 50.930 -8.670 51.460 -8.360 ;
        RECT 52.570 -8.670 52.890 -8.360 ;
        RECT 53.480 -8.670 53.800 -8.360 ;
        RECT 48.960 -9.410 49.280 -9.100 ;
        RECT 49.870 -9.410 50.190 -9.100 ;
        RECT 51.320 -9.190 51.460 -8.670 ;
        RECT 45.180 -11.080 45.710 -10.770 ;
        RECT 46.820 -11.080 47.140 -10.770 ;
        RECT 47.730 -11.080 48.050 -10.770 ;
        RECT 45.570 -12.590 45.710 -11.080 ;
        RECT 45.480 -12.910 45.800 -12.590 ;
        RECT 44.120 -14.570 44.450 -14.240 ;
        RECT 44.210 -19.890 44.350 -14.570 ;
        RECT 44.210 -20.210 44.630 -19.890 ;
        RECT 45.570 -21.780 45.710 -12.910 ;
        RECT 46.190 -14.110 46.510 -13.790 ;
        RECT 46.270 -14.630 46.440 -14.110 ;
        RECT 46.910 -14.240 47.050 -11.080 ;
        RECT 46.830 -14.570 47.160 -14.240 ;
        RECT 46.210 -15.030 46.510 -14.630 ;
        RECT 46.910 -19.890 47.050 -14.570 ;
        RECT 46.620 -20.210 47.050 -19.890 ;
        RECT 45.480 -22.100 45.800 -21.780 ;
        RECT 41.990 -23.030 42.310 -22.710 ;
        RECT 43.210 -23.030 43.530 -22.710 ;
        RECT 33.980 -23.760 34.300 -23.440 ;
        RECT 39.730 -23.760 40.050 -23.440 ;
        RECT 42.550 -23.580 42.950 -23.180 ;
        RECT 45.570 -23.440 45.710 -22.100 ;
        RECT 47.830 -22.710 47.970 -11.080 ;
        RECT 49.050 -22.710 49.190 -9.410 ;
        RECT 49.960 -14.240 50.100 -9.410 ;
        RECT 51.320 -9.500 51.830 -9.190 ;
        RECT 51.320 -10.770 51.460 -9.500 ;
        RECT 52.660 -10.770 52.800 -8.670 ;
        RECT 53.580 -10.770 53.720 -8.670 ;
        RECT 54.800 -9.100 54.940 -7.000 ;
        RECT 55.710 -9.100 55.850 -7.000 ;
        RECT 57.070 -7.090 57.580 -6.780 ;
        RECT 57.070 -8.360 57.210 -7.090 ;
        RECT 58.410 -8.360 58.550 -5.670 ;
        RECT 59.330 -8.360 59.470 -5.670 ;
        RECT 60.550 -6.690 60.690 -4.000 ;
        RECT 61.460 -6.690 61.600 -4.000 ;
        RECT 62.820 -4.090 63.330 -3.780 ;
        RECT 62.820 -5.360 62.960 -4.090 ;
        RECT 64.160 -5.360 64.300 -3.260 ;
        RECT 65.080 -5.360 65.220 -3.260 ;
        RECT 66.300 -3.690 66.440 -1.590 ;
        RECT 67.210 -3.690 67.350 -1.590 ;
        RECT 68.570 -1.680 69.080 -1.370 ;
        RECT 68.570 -2.950 68.710 -1.680 ;
        RECT 69.910 -2.950 70.050 -0.850 ;
        RECT 70.830 -2.950 70.970 -0.850 ;
        RECT 72.050 -1.280 72.190 0.820 ;
        RECT 72.960 -1.280 73.100 0.820 ;
        RECT 74.320 0.730 74.830 1.040 ;
        RECT 74.320 -0.540 74.460 0.730 ;
        RECT 75.660 -0.540 75.800 1.560 ;
        RECT 76.580 -0.540 76.720 1.560 ;
        RECT 77.800 1.130 77.940 3.230 ;
        RECT 78.710 1.130 78.850 3.230 ;
        RECT 80.070 3.140 80.580 3.450 ;
        RECT 80.070 1.870 80.210 3.140 ;
        RECT 81.410 1.870 81.550 3.970 ;
        RECT 82.330 1.870 82.470 3.970 ;
        RECT 83.550 3.540 83.690 5.640 ;
        RECT 84.460 3.540 84.600 5.640 ;
        RECT 85.820 5.550 86.330 5.860 ;
        RECT 85.820 4.280 85.960 5.550 ;
        RECT 87.160 4.280 87.300 6.380 ;
        RECT 88.080 4.280 88.220 6.380 ;
        RECT 89.300 5.950 89.440 8.050 ;
        RECT 90.210 5.950 90.350 8.050 ;
        RECT 91.570 7.960 92.080 8.270 ;
        RECT 91.570 6.690 91.710 7.960 ;
        RECT 92.910 6.690 93.050 9.200 ;
        RECT 93.830 6.690 93.970 9.200 ;
        RECT 91.180 6.380 91.710 6.690 ;
        RECT 92.820 6.380 93.140 6.690 ;
        RECT 93.730 6.380 94.050 6.690 ;
        RECT 89.210 5.640 89.530 5.950 ;
        RECT 90.120 5.640 90.440 5.950 ;
        RECT 91.570 5.860 91.710 6.380 ;
        RECT 85.430 3.970 85.960 4.280 ;
        RECT 87.070 3.970 87.390 4.280 ;
        RECT 87.980 3.970 88.300 4.280 ;
        RECT 83.460 3.230 83.780 3.540 ;
        RECT 84.370 3.230 84.690 3.540 ;
        RECT 85.820 3.450 85.960 3.970 ;
        RECT 79.680 1.560 80.210 1.870 ;
        RECT 81.320 1.560 81.640 1.870 ;
        RECT 82.230 1.560 82.550 1.870 ;
        RECT 77.710 0.820 78.030 1.130 ;
        RECT 78.620 0.820 78.940 1.130 ;
        RECT 80.070 1.040 80.210 1.560 ;
        RECT 73.930 -0.850 74.460 -0.540 ;
        RECT 75.570 -0.850 75.890 -0.540 ;
        RECT 76.480 -0.850 76.800 -0.540 ;
        RECT 71.960 -1.590 72.280 -1.280 ;
        RECT 72.870 -1.590 73.190 -1.280 ;
        RECT 74.320 -1.370 74.460 -0.850 ;
        RECT 68.180 -3.260 68.710 -2.950 ;
        RECT 69.820 -3.260 70.140 -2.950 ;
        RECT 70.730 -3.260 71.050 -2.950 ;
        RECT 66.210 -4.000 66.530 -3.690 ;
        RECT 67.120 -4.000 67.440 -3.690 ;
        RECT 68.570 -3.780 68.710 -3.260 ;
        RECT 62.430 -5.670 62.960 -5.360 ;
        RECT 64.070 -5.670 64.390 -5.360 ;
        RECT 64.980 -5.670 65.300 -5.360 ;
        RECT 60.460 -7.000 60.780 -6.690 ;
        RECT 61.370 -7.000 61.690 -6.690 ;
        RECT 62.820 -6.780 62.960 -5.670 ;
        RECT 56.680 -8.670 57.210 -8.360 ;
        RECT 58.320 -8.670 58.640 -8.360 ;
        RECT 59.230 -8.670 59.550 -8.360 ;
        RECT 54.710 -9.410 55.030 -9.100 ;
        RECT 55.620 -9.410 55.940 -9.100 ;
        RECT 57.070 -9.190 57.210 -8.670 ;
        RECT 50.930 -11.080 51.460 -10.770 ;
        RECT 52.570 -11.080 52.890 -10.770 ;
        RECT 53.480 -11.080 53.800 -10.770 ;
        RECT 51.320 -12.590 51.460 -11.080 ;
        RECT 51.230 -12.910 51.550 -12.590 ;
        RECT 49.870 -14.570 50.200 -14.240 ;
        RECT 49.960 -19.890 50.100 -14.570 ;
        RECT 49.960 -20.210 50.380 -19.890 ;
        RECT 51.320 -21.780 51.460 -12.910 ;
        RECT 51.940 -14.160 52.260 -13.840 ;
        RECT 52.020 -15.460 52.190 -14.160 ;
        RECT 52.660 -14.240 52.800 -11.080 ;
        RECT 52.580 -14.570 52.910 -14.240 ;
        RECT 51.960 -15.860 52.260 -15.460 ;
        RECT 52.660 -19.890 52.800 -14.570 ;
        RECT 52.370 -20.210 52.800 -19.890 ;
        RECT 51.230 -22.100 51.550 -21.780 ;
        RECT 47.740 -23.030 48.060 -22.710 ;
        RECT 48.960 -23.030 49.280 -22.710 ;
        RECT 51.320 -23.440 51.460 -22.100 ;
        RECT 53.580 -22.710 53.720 -11.080 ;
        RECT 54.800 -22.710 54.940 -9.410 ;
        RECT 55.710 -14.240 55.850 -9.410 ;
        RECT 57.070 -9.500 57.580 -9.190 ;
        RECT 57.070 -10.770 57.210 -9.500 ;
        RECT 58.410 -10.770 58.550 -8.670 ;
        RECT 59.330 -10.770 59.470 -8.670 ;
        RECT 60.550 -9.100 60.690 -7.000 ;
        RECT 61.460 -9.100 61.600 -7.000 ;
        RECT 62.820 -7.090 63.330 -6.780 ;
        RECT 62.820 -8.360 62.960 -7.090 ;
        RECT 64.160 -8.360 64.300 -5.670 ;
        RECT 65.080 -8.360 65.220 -5.670 ;
        RECT 66.300 -6.690 66.440 -4.000 ;
        RECT 67.210 -6.690 67.350 -4.000 ;
        RECT 68.570 -4.090 69.080 -3.780 ;
        RECT 68.570 -5.360 68.710 -4.090 ;
        RECT 69.910 -5.360 70.050 -3.260 ;
        RECT 70.830 -5.360 70.970 -3.260 ;
        RECT 72.050 -3.690 72.190 -1.590 ;
        RECT 72.960 -3.690 73.100 -1.590 ;
        RECT 74.320 -1.680 74.830 -1.370 ;
        RECT 74.320 -2.950 74.460 -1.680 ;
        RECT 75.660 -2.950 75.800 -0.850 ;
        RECT 76.580 -2.950 76.720 -0.850 ;
        RECT 77.800 -1.280 77.940 0.820 ;
        RECT 78.710 -1.280 78.850 0.820 ;
        RECT 80.070 0.730 80.580 1.040 ;
        RECT 80.070 -0.540 80.210 0.730 ;
        RECT 81.410 -0.540 81.550 1.560 ;
        RECT 82.330 -0.540 82.470 1.560 ;
        RECT 83.550 1.130 83.690 3.230 ;
        RECT 84.460 1.130 84.600 3.230 ;
        RECT 85.820 3.140 86.330 3.450 ;
        RECT 85.820 1.870 85.960 3.140 ;
        RECT 87.160 1.870 87.300 3.970 ;
        RECT 88.080 1.870 88.220 3.970 ;
        RECT 89.300 3.540 89.440 5.640 ;
        RECT 90.210 3.540 90.350 5.640 ;
        RECT 91.570 5.550 92.080 5.860 ;
        RECT 91.570 4.280 91.710 5.550 ;
        RECT 92.910 4.280 93.050 6.380 ;
        RECT 93.830 4.280 93.970 6.380 ;
        RECT 91.180 3.970 91.710 4.280 ;
        RECT 92.820 3.970 93.140 4.280 ;
        RECT 93.730 3.970 94.050 4.280 ;
        RECT 89.210 3.230 89.530 3.540 ;
        RECT 90.120 3.230 90.440 3.540 ;
        RECT 91.570 3.450 91.710 3.970 ;
        RECT 85.430 1.560 85.960 1.870 ;
        RECT 87.070 1.560 87.390 1.870 ;
        RECT 87.980 1.560 88.300 1.870 ;
        RECT 83.460 0.820 83.780 1.130 ;
        RECT 84.370 0.820 84.690 1.130 ;
        RECT 85.820 1.040 85.960 1.560 ;
        RECT 79.680 -0.850 80.210 -0.540 ;
        RECT 81.320 -0.850 81.640 -0.540 ;
        RECT 82.230 -0.850 82.550 -0.540 ;
        RECT 77.710 -1.590 78.030 -1.280 ;
        RECT 78.620 -1.590 78.940 -1.280 ;
        RECT 80.070 -1.370 80.210 -0.850 ;
        RECT 73.930 -3.260 74.460 -2.950 ;
        RECT 75.570 -3.260 75.890 -2.950 ;
        RECT 76.480 -3.260 76.800 -2.950 ;
        RECT 71.960 -4.000 72.280 -3.690 ;
        RECT 72.870 -4.000 73.190 -3.690 ;
        RECT 74.320 -3.780 74.460 -3.260 ;
        RECT 68.180 -5.670 68.710 -5.360 ;
        RECT 69.820 -5.670 70.140 -5.360 ;
        RECT 70.730 -5.670 71.050 -5.360 ;
        RECT 66.210 -7.000 66.530 -6.690 ;
        RECT 67.120 -7.000 67.440 -6.690 ;
        RECT 68.570 -6.780 68.710 -5.670 ;
        RECT 62.430 -8.670 62.960 -8.360 ;
        RECT 64.070 -8.670 64.390 -8.360 ;
        RECT 64.980 -8.670 65.300 -8.360 ;
        RECT 60.460 -9.410 60.780 -9.100 ;
        RECT 61.370 -9.410 61.690 -9.100 ;
        RECT 62.820 -9.190 62.960 -8.670 ;
        RECT 56.680 -11.080 57.210 -10.770 ;
        RECT 58.320 -11.080 58.640 -10.770 ;
        RECT 59.230 -11.080 59.550 -10.770 ;
        RECT 57.070 -12.590 57.210 -11.080 ;
        RECT 56.980 -12.910 57.300 -12.590 ;
        RECT 55.620 -14.570 55.950 -14.240 ;
        RECT 55.710 -19.890 55.850 -14.570 ;
        RECT 55.710 -20.210 56.130 -19.890 ;
        RECT 57.070 -21.780 57.210 -12.910 ;
        RECT 57.690 -14.130 58.010 -13.810 ;
        RECT 57.770 -16.240 57.940 -14.130 ;
        RECT 58.410 -14.240 58.550 -11.080 ;
        RECT 58.330 -14.570 58.660 -14.240 ;
        RECT 57.710 -16.640 58.010 -16.240 ;
        RECT 58.410 -19.890 58.550 -14.570 ;
        RECT 58.120 -20.210 58.550 -19.890 ;
        RECT 56.980 -22.100 57.300 -21.780 ;
        RECT 53.490 -23.030 53.810 -22.710 ;
        RECT 54.710 -23.030 55.030 -22.710 ;
        RECT 45.480 -23.760 45.800 -23.440 ;
        RECT 51.230 -23.760 51.550 -23.440 ;
        RECT 53.950 -23.560 54.350 -23.160 ;
        RECT 57.070 -23.440 57.210 -22.100 ;
        RECT 59.330 -22.710 59.470 -11.080 ;
        RECT 60.550 -22.710 60.690 -9.410 ;
        RECT 61.460 -14.240 61.600 -9.410 ;
        RECT 62.820 -9.500 63.330 -9.190 ;
        RECT 62.820 -10.770 62.960 -9.500 ;
        RECT 64.160 -10.770 64.300 -8.670 ;
        RECT 65.080 -10.770 65.220 -8.670 ;
        RECT 66.300 -9.100 66.440 -7.000 ;
        RECT 67.210 -9.100 67.350 -7.000 ;
        RECT 68.570 -7.090 69.080 -6.780 ;
        RECT 68.570 -8.360 68.710 -7.090 ;
        RECT 69.910 -8.360 70.050 -5.670 ;
        RECT 70.830 -8.360 70.970 -5.670 ;
        RECT 72.050 -6.690 72.190 -4.000 ;
        RECT 72.960 -6.690 73.100 -4.000 ;
        RECT 74.320 -4.090 74.830 -3.780 ;
        RECT 74.320 -5.360 74.460 -4.090 ;
        RECT 75.660 -5.360 75.800 -3.260 ;
        RECT 76.580 -5.360 76.720 -3.260 ;
        RECT 77.800 -3.690 77.940 -1.590 ;
        RECT 78.710 -3.690 78.850 -1.590 ;
        RECT 80.070 -1.680 80.580 -1.370 ;
        RECT 80.070 -2.950 80.210 -1.680 ;
        RECT 81.410 -2.950 81.550 -0.850 ;
        RECT 82.330 -2.950 82.470 -0.850 ;
        RECT 83.550 -1.280 83.690 0.820 ;
        RECT 84.460 -1.280 84.600 0.820 ;
        RECT 85.820 0.730 86.330 1.040 ;
        RECT 85.820 -0.540 85.960 0.730 ;
        RECT 87.160 -0.540 87.300 1.560 ;
        RECT 88.080 -0.540 88.220 1.560 ;
        RECT 89.300 1.130 89.440 3.230 ;
        RECT 90.210 1.130 90.350 3.230 ;
        RECT 91.570 3.140 92.080 3.450 ;
        RECT 91.570 1.870 91.710 3.140 ;
        RECT 92.910 1.870 93.050 3.970 ;
        RECT 93.830 1.870 93.970 3.970 ;
        RECT 91.180 1.560 91.710 1.870 ;
        RECT 92.820 1.560 93.140 1.870 ;
        RECT 93.730 1.560 94.050 1.870 ;
        RECT 89.210 0.820 89.530 1.130 ;
        RECT 90.120 0.820 90.440 1.130 ;
        RECT 91.570 1.040 91.710 1.560 ;
        RECT 85.430 -0.850 85.960 -0.540 ;
        RECT 87.070 -0.850 87.390 -0.540 ;
        RECT 87.980 -0.850 88.300 -0.540 ;
        RECT 83.460 -1.590 83.780 -1.280 ;
        RECT 84.370 -1.590 84.690 -1.280 ;
        RECT 85.820 -1.370 85.960 -0.850 ;
        RECT 79.680 -3.260 80.210 -2.950 ;
        RECT 81.320 -3.260 81.640 -2.950 ;
        RECT 82.230 -3.260 82.550 -2.950 ;
        RECT 77.710 -4.000 78.030 -3.690 ;
        RECT 78.620 -4.000 78.940 -3.690 ;
        RECT 80.070 -3.780 80.210 -3.260 ;
        RECT 73.930 -5.670 74.460 -5.360 ;
        RECT 75.570 -5.670 75.890 -5.360 ;
        RECT 76.480 -5.670 76.800 -5.360 ;
        RECT 71.960 -7.000 72.280 -6.690 ;
        RECT 72.870 -7.000 73.190 -6.690 ;
        RECT 74.320 -6.780 74.460 -5.670 ;
        RECT 68.180 -8.670 68.710 -8.360 ;
        RECT 69.820 -8.670 70.140 -8.360 ;
        RECT 70.730 -8.670 71.050 -8.360 ;
        RECT 66.210 -9.410 66.530 -9.100 ;
        RECT 67.120 -9.410 67.440 -9.100 ;
        RECT 68.570 -9.190 68.710 -8.670 ;
        RECT 62.430 -11.080 62.960 -10.770 ;
        RECT 64.070 -11.080 64.390 -10.770 ;
        RECT 64.980 -11.080 65.300 -10.770 ;
        RECT 62.820 -12.590 62.960 -11.080 ;
        RECT 62.730 -12.910 63.050 -12.590 ;
        RECT 61.370 -14.570 61.700 -14.240 ;
        RECT 61.460 -19.890 61.600 -14.570 ;
        RECT 61.460 -20.210 61.880 -19.890 ;
        RECT 62.820 -21.780 62.960 -12.910 ;
        RECT 63.440 -14.170 63.760 -13.850 ;
        RECT 63.520 -17.100 63.690 -14.170 ;
        RECT 64.160 -14.240 64.300 -11.080 ;
        RECT 64.080 -14.570 64.410 -14.240 ;
        RECT 63.460 -17.500 63.760 -17.100 ;
        RECT 64.160 -19.890 64.300 -14.570 ;
        RECT 63.870 -20.210 64.300 -19.890 ;
        RECT 62.730 -22.100 63.050 -21.780 ;
        RECT 59.240 -23.030 59.560 -22.710 ;
        RECT 60.460 -23.030 60.780 -22.710 ;
        RECT 62.820 -23.440 62.960 -22.100 ;
        RECT 65.080 -22.710 65.220 -11.080 ;
        RECT 66.300 -22.710 66.440 -9.410 ;
        RECT 67.210 -14.240 67.350 -9.410 ;
        RECT 68.570 -9.500 69.080 -9.190 ;
        RECT 68.570 -10.770 68.710 -9.500 ;
        RECT 69.910 -10.770 70.050 -8.670 ;
        RECT 70.830 -10.770 70.970 -8.670 ;
        RECT 72.050 -9.100 72.190 -7.000 ;
        RECT 72.960 -9.100 73.100 -7.000 ;
        RECT 74.320 -7.090 74.830 -6.780 ;
        RECT 74.320 -8.360 74.460 -7.090 ;
        RECT 75.660 -8.360 75.800 -5.670 ;
        RECT 76.580 -8.360 76.720 -5.670 ;
        RECT 77.800 -6.690 77.940 -4.000 ;
        RECT 78.710 -6.690 78.850 -4.000 ;
        RECT 80.070 -4.090 80.580 -3.780 ;
        RECT 80.070 -5.360 80.210 -4.090 ;
        RECT 81.410 -5.360 81.550 -3.260 ;
        RECT 82.330 -5.360 82.470 -3.260 ;
        RECT 83.550 -3.690 83.690 -1.590 ;
        RECT 84.460 -3.690 84.600 -1.590 ;
        RECT 85.820 -1.680 86.330 -1.370 ;
        RECT 85.820 -2.950 85.960 -1.680 ;
        RECT 87.160 -2.950 87.300 -0.850 ;
        RECT 88.080 -2.950 88.220 -0.850 ;
        RECT 89.300 -1.280 89.440 0.820 ;
        RECT 90.210 -1.280 90.350 0.820 ;
        RECT 91.570 0.730 92.080 1.040 ;
        RECT 91.570 -0.540 91.710 0.730 ;
        RECT 92.910 -0.540 93.050 1.560 ;
        RECT 93.830 -0.540 93.970 1.560 ;
        RECT 91.180 -0.850 91.710 -0.540 ;
        RECT 92.820 -0.850 93.140 -0.540 ;
        RECT 93.730 -0.850 94.050 -0.540 ;
        RECT 89.210 -1.590 89.530 -1.280 ;
        RECT 90.120 -1.590 90.440 -1.280 ;
        RECT 91.570 -1.370 91.710 -0.850 ;
        RECT 85.430 -3.260 85.960 -2.950 ;
        RECT 87.070 -3.260 87.390 -2.950 ;
        RECT 87.980 -3.260 88.300 -2.950 ;
        RECT 83.460 -4.000 83.780 -3.690 ;
        RECT 84.370 -4.000 84.690 -3.690 ;
        RECT 85.820 -3.780 85.960 -3.260 ;
        RECT 79.680 -5.670 80.210 -5.360 ;
        RECT 81.320 -5.670 81.640 -5.360 ;
        RECT 82.230 -5.670 82.550 -5.360 ;
        RECT 77.710 -7.000 78.030 -6.690 ;
        RECT 78.620 -7.000 78.940 -6.690 ;
        RECT 80.070 -6.780 80.210 -5.670 ;
        RECT 73.930 -8.670 74.460 -8.360 ;
        RECT 75.570 -8.670 75.890 -8.360 ;
        RECT 76.480 -8.670 76.800 -8.360 ;
        RECT 71.960 -9.410 72.280 -9.100 ;
        RECT 72.870 -9.410 73.190 -9.100 ;
        RECT 74.320 -9.190 74.460 -8.670 ;
        RECT 68.180 -11.080 68.710 -10.770 ;
        RECT 69.820 -11.080 70.140 -10.770 ;
        RECT 70.730 -11.080 71.050 -10.770 ;
        RECT 68.570 -12.590 68.710 -11.080 ;
        RECT 68.480 -12.910 68.800 -12.590 ;
        RECT 67.120 -14.570 67.450 -14.240 ;
        RECT 67.210 -19.890 67.350 -14.570 ;
        RECT 67.210 -20.210 67.630 -19.890 ;
        RECT 68.570 -21.780 68.710 -12.910 ;
        RECT 69.190 -14.180 69.510 -13.860 ;
        RECT 69.270 -17.900 69.440 -14.180 ;
        RECT 69.910 -14.240 70.050 -11.080 ;
        RECT 69.830 -14.570 70.160 -14.240 ;
        RECT 69.210 -18.300 69.510 -17.900 ;
        RECT 69.910 -19.890 70.050 -14.570 ;
        RECT 69.620 -20.210 70.050 -19.890 ;
        RECT 68.480 -22.100 68.800 -21.780 ;
        RECT 64.990 -23.030 65.310 -22.710 ;
        RECT 66.210 -23.030 66.530 -22.710 ;
        RECT 56.980 -23.760 57.300 -23.440 ;
        RECT 62.730 -23.760 63.050 -23.440 ;
        RECT 65.630 -23.560 66.030 -23.160 ;
        RECT 68.570 -23.440 68.710 -22.100 ;
        RECT 70.830 -22.710 70.970 -11.080 ;
        RECT 72.050 -22.710 72.190 -9.410 ;
        RECT 72.960 -14.240 73.100 -9.410 ;
        RECT 74.320 -9.500 74.830 -9.190 ;
        RECT 74.320 -10.770 74.460 -9.500 ;
        RECT 75.660 -10.770 75.800 -8.670 ;
        RECT 76.580 -10.770 76.720 -8.670 ;
        RECT 77.800 -9.100 77.940 -7.000 ;
        RECT 78.710 -9.100 78.850 -7.000 ;
        RECT 80.070 -7.090 80.580 -6.780 ;
        RECT 80.070 -8.360 80.210 -7.090 ;
        RECT 81.410 -8.360 81.550 -5.670 ;
        RECT 82.330 -8.360 82.470 -5.670 ;
        RECT 83.550 -6.690 83.690 -4.000 ;
        RECT 84.460 -6.690 84.600 -4.000 ;
        RECT 85.820 -4.090 86.330 -3.780 ;
        RECT 85.820 -5.360 85.960 -4.090 ;
        RECT 87.160 -5.360 87.300 -3.260 ;
        RECT 88.080 -5.360 88.220 -3.260 ;
        RECT 89.300 -3.690 89.440 -1.590 ;
        RECT 90.210 -3.690 90.350 -1.590 ;
        RECT 91.570 -1.680 92.080 -1.370 ;
        RECT 91.570 -2.950 91.710 -1.680 ;
        RECT 92.910 -2.950 93.050 -0.850 ;
        RECT 93.830 -2.950 93.970 -0.850 ;
        RECT 91.180 -3.260 91.710 -2.950 ;
        RECT 92.820 -3.260 93.140 -2.950 ;
        RECT 93.730 -3.260 94.050 -2.950 ;
        RECT 89.210 -4.000 89.530 -3.690 ;
        RECT 90.120 -4.000 90.440 -3.690 ;
        RECT 91.570 -3.780 91.710 -3.260 ;
        RECT 85.430 -5.670 85.960 -5.360 ;
        RECT 87.070 -5.670 87.390 -5.360 ;
        RECT 87.980 -5.670 88.300 -5.360 ;
        RECT 83.460 -7.000 83.780 -6.690 ;
        RECT 84.370 -7.000 84.690 -6.690 ;
        RECT 85.820 -6.780 85.960 -5.670 ;
        RECT 79.680 -8.670 80.210 -8.360 ;
        RECT 81.320 -8.670 81.640 -8.360 ;
        RECT 82.230 -8.670 82.550 -8.360 ;
        RECT 77.710 -9.410 78.030 -9.100 ;
        RECT 78.620 -9.410 78.940 -9.100 ;
        RECT 80.070 -9.190 80.210 -8.670 ;
        RECT 73.930 -11.080 74.460 -10.770 ;
        RECT 75.570 -11.080 75.890 -10.770 ;
        RECT 76.480 -11.080 76.800 -10.770 ;
        RECT 74.320 -12.590 74.460 -11.080 ;
        RECT 74.230 -12.910 74.550 -12.590 ;
        RECT 72.870 -14.570 73.200 -14.240 ;
        RECT 72.960 -19.890 73.100 -14.570 ;
        RECT 72.960 -20.210 73.380 -19.890 ;
        RECT 74.320 -21.780 74.460 -12.910 ;
        RECT 74.940 -14.140 75.260 -13.820 ;
        RECT 75.020 -18.700 75.190 -14.140 ;
        RECT 75.660 -14.240 75.800 -11.080 ;
        RECT 75.580 -14.570 75.910 -14.240 ;
        RECT 74.960 -19.100 75.260 -18.700 ;
        RECT 75.660 -19.890 75.800 -14.570 ;
        RECT 75.370 -20.210 75.800 -19.890 ;
        RECT 74.230 -22.100 74.550 -21.780 ;
        RECT 70.740 -23.030 71.060 -22.710 ;
        RECT 71.960 -23.030 72.280 -22.710 ;
        RECT 74.320 -23.440 74.460 -22.100 ;
        RECT 76.580 -22.710 76.720 -11.080 ;
        RECT 77.800 -22.710 77.940 -9.410 ;
        RECT 78.710 -14.240 78.850 -9.410 ;
        RECT 80.070 -9.500 80.580 -9.190 ;
        RECT 80.070 -10.770 80.210 -9.500 ;
        RECT 81.410 -10.770 81.550 -8.670 ;
        RECT 82.330 -10.770 82.470 -8.670 ;
        RECT 83.550 -9.100 83.690 -7.000 ;
        RECT 84.460 -9.100 84.600 -7.000 ;
        RECT 85.820 -7.090 86.330 -6.780 ;
        RECT 85.820 -8.360 85.960 -7.090 ;
        RECT 87.160 -8.360 87.300 -5.670 ;
        RECT 88.080 -8.360 88.220 -5.670 ;
        RECT 89.300 -6.690 89.440 -4.000 ;
        RECT 90.210 -6.690 90.350 -4.000 ;
        RECT 91.570 -4.090 92.080 -3.780 ;
        RECT 91.570 -5.360 91.710 -4.090 ;
        RECT 92.910 -5.360 93.050 -3.260 ;
        RECT 93.830 -5.360 93.970 -3.260 ;
        RECT 91.180 -5.670 91.710 -5.360 ;
        RECT 92.820 -5.670 93.140 -5.360 ;
        RECT 93.730 -5.670 94.050 -5.360 ;
        RECT 89.210 -7.000 89.530 -6.690 ;
        RECT 90.120 -7.000 90.440 -6.690 ;
        RECT 91.570 -6.780 91.710 -5.670 ;
        RECT 85.430 -8.670 85.960 -8.360 ;
        RECT 87.070 -8.670 87.390 -8.360 ;
        RECT 87.980 -8.670 88.300 -8.360 ;
        RECT 83.460 -9.410 83.780 -9.100 ;
        RECT 84.370 -9.410 84.690 -9.100 ;
        RECT 85.820 -9.190 85.960 -8.670 ;
        RECT 79.680 -11.080 80.210 -10.770 ;
        RECT 81.320 -11.080 81.640 -10.770 ;
        RECT 82.230 -11.080 82.550 -10.770 ;
        RECT 80.070 -12.590 80.210 -11.080 ;
        RECT 79.980 -12.910 80.300 -12.590 ;
        RECT 78.620 -14.570 78.950 -14.240 ;
        RECT 78.710 -19.890 78.850 -14.570 ;
        RECT 78.710 -20.210 79.130 -19.890 ;
        RECT 80.070 -21.780 80.210 -12.910 ;
        RECT 80.690 -14.180 81.010 -13.860 ;
        RECT 80.770 -19.350 80.940 -14.180 ;
        RECT 81.410 -14.240 81.550 -11.080 ;
        RECT 81.330 -14.570 81.660 -14.240 ;
        RECT 80.710 -19.750 81.010 -19.350 ;
        RECT 81.410 -19.890 81.550 -14.570 ;
        RECT 81.120 -20.210 81.550 -19.890 ;
        RECT 79.980 -22.100 80.300 -21.780 ;
        RECT 76.490 -23.030 76.810 -22.710 ;
        RECT 77.710 -23.030 78.030 -22.710 ;
        RECT 68.480 -23.760 68.800 -23.440 ;
        RECT 74.230 -23.760 74.550 -23.440 ;
        RECT 77.080 -23.560 77.480 -23.160 ;
        RECT 80.070 -23.440 80.210 -22.100 ;
        RECT 82.330 -22.710 82.470 -11.080 ;
        RECT 83.550 -22.710 83.690 -9.410 ;
        RECT 84.460 -14.240 84.600 -9.410 ;
        RECT 85.820 -9.500 86.330 -9.190 ;
        RECT 85.820 -10.770 85.960 -9.500 ;
        RECT 87.160 -10.770 87.300 -8.670 ;
        RECT 88.080 -10.770 88.220 -8.670 ;
        RECT 89.300 -9.100 89.440 -7.000 ;
        RECT 90.210 -9.100 90.350 -7.000 ;
        RECT 91.570 -7.090 92.080 -6.780 ;
        RECT 91.570 -8.360 91.710 -7.090 ;
        RECT 92.910 -8.360 93.050 -5.670 ;
        RECT 93.830 -8.360 93.970 -5.670 ;
        RECT 91.180 -8.670 91.710 -8.360 ;
        RECT 92.820 -8.670 93.140 -8.360 ;
        RECT 93.730 -8.670 94.050 -8.360 ;
        RECT 89.210 -9.410 89.530 -9.100 ;
        RECT 90.120 -9.410 90.440 -9.100 ;
        RECT 91.570 -9.190 91.710 -8.670 ;
        RECT 85.430 -11.080 85.960 -10.770 ;
        RECT 87.070 -11.080 87.390 -10.770 ;
        RECT 87.980 -11.080 88.300 -10.770 ;
        RECT 85.820 -12.590 85.960 -11.080 ;
        RECT 85.730 -12.910 86.050 -12.590 ;
        RECT 84.370 -14.570 84.700 -14.240 ;
        RECT 84.460 -19.890 84.600 -14.570 ;
        RECT 84.460 -20.210 84.880 -19.890 ;
        RECT 85.820 -21.780 85.960 -12.910 ;
        RECT 86.440 -14.140 86.760 -13.820 ;
        RECT 86.520 -20.490 86.690 -14.140 ;
        RECT 87.160 -14.240 87.300 -11.080 ;
        RECT 87.080 -14.570 87.410 -14.240 ;
        RECT 87.160 -19.890 87.300 -14.570 ;
        RECT 86.870 -20.210 87.300 -19.890 ;
        RECT 86.460 -20.890 86.760 -20.490 ;
        RECT 85.730 -22.100 86.050 -21.780 ;
        RECT 82.240 -23.030 82.560 -22.710 ;
        RECT 83.460 -23.030 83.780 -22.710 ;
        RECT 85.820 -23.440 85.960 -22.100 ;
        RECT 88.080 -22.710 88.220 -11.080 ;
        RECT 89.300 -22.710 89.440 -9.410 ;
        RECT 90.210 -14.240 90.350 -9.410 ;
        RECT 91.570 -9.500 92.080 -9.190 ;
        RECT 91.570 -10.770 91.710 -9.500 ;
        RECT 92.910 -10.770 93.050 -8.670 ;
        RECT 93.830 -10.770 93.970 -8.670 ;
        RECT 91.180 -11.080 91.710 -10.770 ;
        RECT 92.820 -11.080 93.140 -10.770 ;
        RECT 93.730 -11.080 94.050 -10.770 ;
        RECT 91.570 -12.590 91.710 -11.080 ;
        RECT 91.480 -12.910 91.800 -12.590 ;
        RECT 90.120 -14.570 90.450 -14.240 ;
        RECT 90.210 -19.890 90.350 -14.570 ;
        RECT 90.210 -20.210 90.630 -19.890 ;
        RECT 91.570 -21.780 91.710 -12.910 ;
        RECT 92.190 -14.150 92.510 -13.830 ;
        RECT 92.270 -21.380 92.440 -14.150 ;
        RECT 92.910 -14.240 93.050 -11.080 ;
        RECT 92.830 -14.570 93.160 -14.240 ;
        RECT 92.910 -19.890 93.050 -14.570 ;
        RECT 92.620 -20.210 93.050 -19.890 ;
        RECT 92.210 -21.780 92.510 -21.380 ;
        RECT 91.480 -22.100 91.800 -21.780 ;
        RECT 87.990 -23.030 88.310 -22.710 ;
        RECT 89.210 -23.030 89.530 -22.710 ;
        RECT 79.980 -23.760 80.300 -23.440 ;
        RECT 85.730 -23.760 86.050 -23.440 ;
        RECT 88.650 -23.540 89.050 -23.140 ;
        RECT 91.570 -23.440 91.710 -22.100 ;
        RECT 93.830 -22.710 93.970 -11.080 ;
        RECT 93.740 -23.030 94.060 -22.710 ;
        RECT 91.480 -23.760 91.800 -23.440 ;
        RECT 7.300 -24.540 7.700 -24.140 ;
        RECT 8.850 -24.540 9.250 -24.140 ;
        RECT 18.800 -24.540 19.200 -24.140 ;
        RECT 20.350 -24.540 20.750 -24.140 ;
        RECT 30.300 -24.540 30.700 -24.140 ;
        RECT 31.840 -24.540 32.240 -24.140 ;
        RECT 41.770 -24.540 42.170 -24.140 ;
        RECT 43.360 -24.550 43.760 -24.150 ;
        RECT 53.290 -24.540 53.690 -24.140 ;
        RECT 54.840 -24.540 55.240 -24.140 ;
        RECT 64.800 -24.550 65.200 -24.150 ;
        RECT 66.330 -24.550 66.730 -24.150 ;
        RECT 76.310 -24.540 76.710 -24.140 ;
        RECT 77.840 -24.540 78.240 -24.140 ;
        RECT 87.800 -24.540 88.200 -24.140 ;
        RECT 89.320 -24.540 89.720 -24.130 ;
        RECT -39.270 -24.870 -38.950 -24.550 ;
        RECT -39.180 -41.280 -39.040 -24.870 ;
        RECT 4.610 -25.310 5.010 -24.910 ;
        RECT 11.540 -25.240 11.940 -24.840 ;
        RECT 16.100 -25.230 16.500 -24.830 ;
        RECT 23.030 -25.280 23.430 -24.880 ;
        RECT 27.620 -25.290 28.020 -24.890 ;
        RECT 34.540 -25.270 34.940 -24.870 ;
        RECT 39.120 -25.290 39.520 -24.890 ;
        RECT 46.030 -25.310 46.430 -24.910 ;
        RECT 50.610 -25.250 51.010 -24.850 ;
        RECT 57.540 -25.270 57.940 -24.870 ;
        RECT 62.110 -25.230 62.510 -24.830 ;
        RECT 69.030 -25.270 69.430 -24.870 ;
        RECT 73.610 -25.270 74.010 -24.870 ;
        RECT 80.530 -25.300 80.930 -24.900 ;
        RECT 85.110 -25.290 85.510 -24.890 ;
        RECT 92.030 -25.250 92.390 -24.870 ;
        RECT -27.470 -25.690 -27.150 -25.370 ;
        RECT 135.320 -25.660 135.580 -25.340 ;
        RECT -35.240 -31.020 -34.940 -30.620 ;
        RECT -35.160 -33.580 -35.020 -31.020 ;
        RECT -35.250 -33.900 -34.930 -33.580 ;
        RECT -39.300 -41.660 -38.920 -41.280 ;
        RECT -41.780 -43.750 -41.520 -43.430 ;
        RECT -39.130 -43.750 -38.870 -43.430 ;
        RECT -39.070 -46.330 -38.930 -43.750 ;
        RECT -37.900 -44.240 -37.580 -43.920 ;
        RECT -39.130 -46.650 -38.870 -46.330 ;
        RECT -39.070 -70.760 -38.930 -46.650 ;
        RECT -37.820 -48.460 -37.680 -44.240 ;
        RECT -37.910 -48.780 -37.590 -48.460 ;
        RECT -37.820 -66.040 -37.680 -48.780 ;
        RECT -35.160 -56.180 -35.020 -33.900 ;
        RECT -27.390 -41.320 -27.220 -25.690 ;
        RECT -15.650 -26.320 -15.390 -26.000 ;
        RECT 125.830 -26.130 126.150 -25.870 ;
        RECT -23.740 -31.020 -23.440 -30.620 ;
        RECT -23.660 -33.580 -23.520 -31.020 ;
        RECT -23.750 -33.900 -23.430 -33.580 ;
        RECT -27.460 -41.640 -27.140 -41.320 ;
        RECT -32.910 -43.750 -32.650 -43.430 ;
        RECT -32.850 -44.930 -32.710 -43.750 ;
        RECT -26.400 -44.240 -26.080 -43.920 ;
        RECT -32.890 -45.250 -32.610 -44.930 ;
        RECT -32.850 -46.360 -32.710 -45.250 ;
        RECT -32.940 -46.620 -32.620 -46.360 ;
        RECT -26.320 -48.460 -26.180 -44.240 ;
        RECT -26.410 -48.780 -26.090 -48.460 ;
        RECT -35.250 -56.500 -34.930 -56.180 ;
        RECT -35.160 -60.910 -35.020 -56.500 ;
        RECT -35.250 -61.230 -34.930 -60.910 ;
        RECT -37.900 -66.360 -37.580 -66.040 ;
        RECT -37.830 -68.630 -37.690 -68.620 ;
        RECT -37.910 -68.950 -37.590 -68.630 ;
        RECT -39.130 -71.080 -38.870 -70.760 ;
        RECT -39.070 -73.690 -38.930 -71.080 ;
        RECT -39.160 -73.950 -38.840 -73.690 ;
        RECT -37.830 -75.800 -37.690 -68.950 ;
        RECT -37.910 -76.120 -37.590 -75.800 ;
        RECT -35.160 -83.510 -35.020 -61.230 ;
        RECT -26.320 -66.040 -26.180 -48.780 ;
        RECT -23.660 -56.180 -23.520 -33.900 ;
        RECT -15.600 -41.320 -15.430 -26.320 ;
        RECT 114.200 -26.630 114.520 -26.370 ;
        RECT -3.870 -27.070 -3.610 -26.750 ;
        RECT -11.840 -33.580 -11.700 -31.170 ;
        RECT -11.930 -33.900 -11.610 -33.580 ;
        RECT -15.640 -41.640 -15.380 -41.320 ;
        RECT -21.410 -43.750 -21.150 -43.430 ;
        RECT -21.350 -44.930 -21.210 -43.750 ;
        RECT -14.580 -44.240 -14.260 -43.920 ;
        RECT -21.390 -45.250 -21.110 -44.930 ;
        RECT -21.350 -46.360 -21.210 -45.250 ;
        RECT -21.440 -46.620 -21.120 -46.360 ;
        RECT -14.500 -48.460 -14.360 -44.240 ;
        RECT -14.590 -48.780 -14.270 -48.460 ;
        RECT -23.750 -56.500 -23.430 -56.180 ;
        RECT -23.660 -60.910 -23.520 -56.500 ;
        RECT -23.750 -61.230 -23.430 -60.910 ;
        RECT -26.400 -66.360 -26.080 -66.040 ;
        RECT -26.330 -68.630 -26.190 -68.620 ;
        RECT -26.410 -68.950 -26.090 -68.630 ;
        RECT -32.970 -71.080 -32.710 -70.760 ;
        RECT -32.910 -72.270 -32.770 -71.080 ;
        RECT -32.910 -72.590 -32.650 -72.270 ;
        RECT -32.910 -73.660 -32.770 -72.590 ;
        RECT -33.000 -73.980 -32.680 -73.660 ;
        RECT -26.330 -75.800 -26.190 -68.950 ;
        RECT -26.410 -76.120 -26.090 -75.800 ;
        RECT -23.660 -83.510 -23.520 -61.230 ;
        RECT -14.500 -66.040 -14.360 -48.780 ;
        RECT -11.840 -56.180 -11.700 -33.900 ;
        RECT -3.820 -41.320 -3.650 -27.070 ;
        RECT 102.070 -27.260 102.390 -27.000 ;
        RECT 8.080 -27.780 8.400 -27.460 ;
        RECT -0.110 -31.060 0.190 -30.660 ;
        RECT -0.030 -33.580 0.110 -31.060 ;
        RECT -0.120 -33.900 0.200 -33.580 ;
        RECT -3.860 -41.640 -3.600 -41.320 ;
        RECT -9.590 -43.750 -9.330 -43.430 ;
        RECT -9.530 -44.930 -9.390 -43.750 ;
        RECT -2.770 -44.240 -2.450 -43.920 ;
        RECT -9.570 -45.250 -9.290 -44.930 ;
        RECT -9.530 -46.360 -9.390 -45.250 ;
        RECT -9.620 -46.620 -9.300 -46.360 ;
        RECT -2.690 -48.460 -2.550 -44.240 ;
        RECT -2.780 -48.780 -2.460 -48.460 ;
        RECT -11.930 -56.500 -11.610 -56.180 ;
        RECT -11.840 -60.910 -11.700 -56.500 ;
        RECT -11.930 -61.230 -11.610 -60.910 ;
        RECT -14.580 -66.360 -14.260 -66.040 ;
        RECT -14.510 -68.630 -14.370 -68.620 ;
        RECT -14.590 -68.950 -14.270 -68.630 ;
        RECT -21.470 -71.080 -21.210 -70.760 ;
        RECT -21.410 -72.270 -21.270 -71.080 ;
        RECT -21.410 -72.590 -21.150 -72.270 ;
        RECT -21.410 -73.660 -21.270 -72.590 ;
        RECT -21.500 -73.980 -21.180 -73.660 ;
        RECT -14.510 -75.800 -14.370 -68.950 ;
        RECT -14.590 -76.120 -14.270 -75.800 ;
        RECT -11.840 -83.510 -11.700 -61.230 ;
        RECT -2.690 -66.040 -2.550 -48.780 ;
        RECT -0.030 -56.180 0.110 -33.900 ;
        RECT 8.160 -41.320 8.330 -27.780 ;
        RECT 90.330 -27.890 90.650 -27.630 ;
        RECT 19.750 -28.580 20.070 -28.260 ;
        RECT 11.700 -31.040 12.000 -30.640 ;
        RECT 11.780 -33.580 11.920 -31.040 ;
        RECT 11.690 -33.900 12.010 -33.580 ;
        RECT 8.090 -41.640 8.410 -41.320 ;
        RECT 2.220 -43.750 2.480 -43.430 ;
        RECT 2.280 -44.930 2.420 -43.750 ;
        RECT 9.040 -44.240 9.360 -43.920 ;
        RECT 2.240 -45.250 2.520 -44.930 ;
        RECT 2.280 -46.360 2.420 -45.250 ;
        RECT 2.190 -46.620 2.510 -46.360 ;
        RECT 9.120 -48.460 9.260 -44.240 ;
        RECT 9.030 -48.780 9.350 -48.460 ;
        RECT -0.120 -56.500 0.200 -56.180 ;
        RECT -0.030 -60.910 0.110 -56.500 ;
        RECT -0.120 -61.230 0.200 -60.910 ;
        RECT -2.770 -66.360 -2.450 -66.040 ;
        RECT -2.700 -68.630 -2.560 -68.620 ;
        RECT -2.780 -68.950 -2.460 -68.630 ;
        RECT -9.650 -71.080 -9.390 -70.760 ;
        RECT -9.590 -72.270 -9.450 -71.080 ;
        RECT -9.590 -72.590 -9.330 -72.270 ;
        RECT -9.590 -73.660 -9.450 -72.590 ;
        RECT -9.680 -73.980 -9.360 -73.660 ;
        RECT -2.700 -75.800 -2.560 -68.950 ;
        RECT -2.780 -76.120 -2.460 -75.800 ;
        RECT -0.030 -83.510 0.110 -61.230 ;
        RECT 9.120 -66.040 9.260 -48.780 ;
        RECT 11.780 -56.180 11.920 -33.900 ;
        RECT 19.830 -41.310 20.000 -28.580 ;
        RECT 78.480 -28.640 78.740 -28.320 ;
        RECT 31.340 -29.420 31.660 -29.100 ;
        RECT 23.520 -31.050 23.820 -30.650 ;
        RECT 23.600 -33.580 23.740 -31.050 ;
        RECT 23.510 -33.900 23.830 -33.580 ;
        RECT 19.750 -41.630 20.080 -41.310 ;
        RECT 14.030 -43.750 14.290 -43.430 ;
        RECT 14.090 -44.930 14.230 -43.750 ;
        RECT 20.860 -44.240 21.180 -43.920 ;
        RECT 14.050 -45.250 14.330 -44.930 ;
        RECT 14.090 -46.360 14.230 -45.250 ;
        RECT 14.000 -46.620 14.320 -46.360 ;
        RECT 20.940 -48.460 21.080 -44.240 ;
        RECT 20.850 -48.780 21.170 -48.460 ;
        RECT 11.690 -56.500 12.010 -56.180 ;
        RECT 11.780 -60.910 11.920 -56.500 ;
        RECT 11.690 -61.230 12.010 -60.910 ;
        RECT 9.040 -66.360 9.360 -66.040 ;
        RECT 9.110 -68.630 9.250 -68.620 ;
        RECT 9.030 -68.950 9.350 -68.630 ;
        RECT 2.160 -71.080 2.420 -70.760 ;
        RECT 2.220 -72.270 2.360 -71.080 ;
        RECT 2.220 -72.590 2.480 -72.270 ;
        RECT 2.220 -73.660 2.360 -72.590 ;
        RECT 2.130 -73.980 2.450 -73.660 ;
        RECT 9.110 -75.800 9.250 -68.950 ;
        RECT 9.030 -76.120 9.350 -75.800 ;
        RECT 11.780 -83.510 11.920 -61.230 ;
        RECT 20.940 -66.040 21.080 -48.780 ;
        RECT 23.600 -56.180 23.740 -33.900 ;
        RECT 31.420 -41.300 31.590 -29.420 ;
        RECT 66.460 -29.440 66.720 -29.120 ;
        RECT 43.080 -30.130 43.400 -29.810 ;
        RECT 35.340 -31.050 35.640 -30.650 ;
        RECT 35.420 -33.580 35.560 -31.050 ;
        RECT 35.330 -33.900 35.650 -33.580 ;
        RECT 31.350 -41.620 31.670 -41.300 ;
        RECT 25.850 -43.750 26.110 -43.430 ;
        RECT 25.910 -44.930 26.050 -43.750 ;
        RECT 32.680 -44.240 33.000 -43.920 ;
        RECT 25.870 -45.250 26.150 -44.930 ;
        RECT 25.910 -46.360 26.050 -45.250 ;
        RECT 25.820 -46.620 26.140 -46.360 ;
        RECT 32.760 -48.460 32.900 -44.240 ;
        RECT 32.670 -48.780 32.990 -48.460 ;
        RECT 23.510 -56.500 23.830 -56.180 ;
        RECT 23.600 -60.910 23.740 -56.500 ;
        RECT 23.510 -61.230 23.830 -60.910 ;
        RECT 20.860 -66.360 21.180 -66.040 ;
        RECT 20.930 -68.630 21.070 -68.620 ;
        RECT 20.850 -68.950 21.170 -68.630 ;
        RECT 13.970 -71.080 14.230 -70.760 ;
        RECT 14.030 -72.270 14.170 -71.080 ;
        RECT 14.030 -72.590 14.290 -72.270 ;
        RECT 14.030 -73.660 14.170 -72.590 ;
        RECT 13.940 -73.980 14.260 -73.660 ;
        RECT 20.930 -75.800 21.070 -68.950 ;
        RECT 20.850 -76.120 21.170 -75.800 ;
        RECT 23.600 -83.510 23.740 -61.230 ;
        RECT 32.760 -66.040 32.900 -48.780 ;
        RECT 35.420 -56.180 35.560 -33.900 ;
        RECT 43.160 -41.300 43.330 -30.130 ;
        RECT 54.960 -30.310 55.220 -29.990 ;
        RECT 47.160 -31.020 47.460 -30.620 ;
        RECT 47.240 -33.580 47.380 -31.020 ;
        RECT 47.150 -33.900 47.470 -33.580 ;
        RECT 43.090 -41.620 43.410 -41.300 ;
        RECT 37.670 -43.750 37.930 -43.430 ;
        RECT 37.730 -44.930 37.870 -43.750 ;
        RECT 44.500 -44.240 44.820 -43.920 ;
        RECT 37.690 -45.250 37.970 -44.930 ;
        RECT 37.730 -46.360 37.870 -45.250 ;
        RECT 37.640 -46.620 37.960 -46.360 ;
        RECT 44.580 -48.460 44.720 -44.240 ;
        RECT 44.490 -48.780 44.810 -48.460 ;
        RECT 35.330 -56.500 35.650 -56.180 ;
        RECT 35.420 -60.910 35.560 -56.500 ;
        RECT 35.330 -61.230 35.650 -60.910 ;
        RECT 32.680 -66.360 33.000 -66.040 ;
        RECT 32.750 -68.630 32.890 -68.620 ;
        RECT 32.670 -68.950 32.990 -68.630 ;
        RECT 25.790 -71.080 26.050 -70.760 ;
        RECT 25.850 -72.270 25.990 -71.080 ;
        RECT 25.850 -72.590 26.110 -72.270 ;
        RECT 25.850 -73.660 25.990 -72.590 ;
        RECT 25.760 -73.980 26.080 -73.660 ;
        RECT 32.750 -75.800 32.890 -68.950 ;
        RECT 32.670 -76.120 32.990 -75.800 ;
        RECT 35.420 -83.510 35.560 -61.230 ;
        RECT 44.580 -66.040 44.720 -48.780 ;
        RECT 47.240 -56.180 47.380 -33.900 ;
        RECT 55.010 -41.300 55.180 -30.310 ;
        RECT 58.980 -31.050 59.280 -30.650 ;
        RECT 59.060 -33.580 59.200 -31.050 ;
        RECT 58.970 -33.900 59.290 -33.580 ;
        RECT 54.970 -41.620 55.230 -41.300 ;
        RECT 49.490 -43.750 49.750 -43.430 ;
        RECT 49.550 -44.930 49.690 -43.750 ;
        RECT 56.320 -44.240 56.640 -43.920 ;
        RECT 49.510 -45.250 49.790 -44.930 ;
        RECT 49.550 -46.360 49.690 -45.250 ;
        RECT 49.460 -46.620 49.780 -46.360 ;
        RECT 56.400 -48.460 56.540 -44.240 ;
        RECT 56.310 -48.780 56.630 -48.460 ;
        RECT 47.150 -56.500 47.470 -56.180 ;
        RECT 47.240 -60.910 47.380 -56.500 ;
        RECT 47.150 -61.230 47.470 -60.910 ;
        RECT 44.500 -66.360 44.820 -66.040 ;
        RECT 44.570 -68.630 44.710 -68.620 ;
        RECT 44.490 -68.950 44.810 -68.630 ;
        RECT 37.610 -71.080 37.870 -70.760 ;
        RECT 37.670 -72.270 37.810 -71.080 ;
        RECT 37.670 -72.590 37.930 -72.270 ;
        RECT 37.670 -73.660 37.810 -72.590 ;
        RECT 37.580 -73.980 37.900 -73.660 ;
        RECT 44.570 -75.800 44.710 -68.950 ;
        RECT 44.490 -76.120 44.810 -75.800 ;
        RECT 47.240 -83.510 47.380 -61.230 ;
        RECT 56.400 -66.040 56.540 -48.780 ;
        RECT 59.060 -56.180 59.200 -33.900 ;
        RECT 66.510 -41.320 66.680 -29.440 ;
        RECT 70.800 -31.050 71.100 -30.650 ;
        RECT 70.880 -33.580 71.020 -31.050 ;
        RECT 70.790 -33.900 71.110 -33.580 ;
        RECT 66.470 -41.640 66.730 -41.320 ;
        RECT 61.310 -43.750 61.570 -43.430 ;
        RECT 61.370 -44.930 61.510 -43.750 ;
        RECT 68.140 -44.240 68.460 -43.920 ;
        RECT 61.330 -45.250 61.610 -44.930 ;
        RECT 61.370 -46.360 61.510 -45.250 ;
        RECT 61.280 -46.620 61.600 -46.360 ;
        RECT 68.220 -48.460 68.360 -44.240 ;
        RECT 68.130 -48.780 68.450 -48.460 ;
        RECT 58.970 -56.500 59.290 -56.180 ;
        RECT 59.060 -60.910 59.200 -56.500 ;
        RECT 58.970 -61.230 59.290 -60.910 ;
        RECT 56.320 -66.360 56.640 -66.040 ;
        RECT 56.390 -68.630 56.530 -68.620 ;
        RECT 56.310 -68.950 56.630 -68.630 ;
        RECT 49.430 -71.080 49.690 -70.760 ;
        RECT 49.490 -72.270 49.630 -71.080 ;
        RECT 49.490 -72.590 49.750 -72.270 ;
        RECT 49.490 -73.660 49.630 -72.590 ;
        RECT 49.400 -73.980 49.720 -73.660 ;
        RECT 56.390 -75.800 56.530 -68.950 ;
        RECT 56.310 -76.120 56.630 -75.800 ;
        RECT 59.060 -83.510 59.200 -61.230 ;
        RECT 68.220 -66.040 68.360 -48.780 ;
        RECT 70.880 -56.180 71.020 -33.900 ;
        RECT 78.530 -41.320 78.700 -28.640 ;
        RECT 82.620 -31.030 82.920 -30.630 ;
        RECT 82.700 -33.580 82.840 -31.030 ;
        RECT 82.610 -33.900 82.930 -33.580 ;
        RECT 78.490 -41.640 78.750 -41.320 ;
        RECT 73.130 -43.750 73.390 -43.430 ;
        RECT 73.190 -44.930 73.330 -43.750 ;
        RECT 79.960 -44.240 80.280 -43.920 ;
        RECT 73.150 -45.250 73.430 -44.930 ;
        RECT 73.190 -46.360 73.330 -45.250 ;
        RECT 73.100 -46.620 73.420 -46.360 ;
        RECT 80.040 -48.460 80.180 -44.240 ;
        RECT 79.950 -48.780 80.270 -48.460 ;
        RECT 70.790 -56.500 71.110 -56.180 ;
        RECT 70.880 -60.910 71.020 -56.500 ;
        RECT 70.790 -61.230 71.110 -60.910 ;
        RECT 68.140 -66.360 68.460 -66.040 ;
        RECT 68.210 -68.630 68.350 -68.620 ;
        RECT 68.130 -68.950 68.450 -68.630 ;
        RECT 61.250 -71.080 61.510 -70.760 ;
        RECT 61.310 -72.270 61.450 -71.080 ;
        RECT 61.310 -72.590 61.570 -72.270 ;
        RECT 61.310 -73.660 61.450 -72.590 ;
        RECT 61.220 -73.980 61.540 -73.660 ;
        RECT 68.210 -75.800 68.350 -68.950 ;
        RECT 68.130 -76.120 68.450 -75.800 ;
        RECT 70.880 -83.510 71.020 -61.230 ;
        RECT 80.040 -66.040 80.180 -48.780 ;
        RECT 82.700 -56.180 82.840 -33.900 ;
        RECT 90.410 -41.350 90.580 -27.890 ;
        RECT 94.460 -31.040 94.760 -30.640 ;
        RECT 94.540 -33.580 94.680 -31.040 ;
        RECT 94.450 -33.900 94.770 -33.580 ;
        RECT 90.340 -41.610 90.660 -41.350 ;
        RECT 84.950 -43.750 85.210 -43.430 ;
        RECT 85.010 -44.930 85.150 -43.750 ;
        RECT 91.800 -44.240 92.120 -43.920 ;
        RECT 84.970 -45.250 85.250 -44.930 ;
        RECT 85.010 -46.360 85.150 -45.250 ;
        RECT 84.920 -46.620 85.240 -46.360 ;
        RECT 91.880 -48.460 92.020 -44.240 ;
        RECT 91.790 -48.780 92.110 -48.460 ;
        RECT 82.610 -56.500 82.930 -56.180 ;
        RECT 82.700 -60.910 82.840 -56.500 ;
        RECT 82.610 -61.230 82.930 -60.910 ;
        RECT 79.960 -66.360 80.280 -66.040 ;
        RECT 80.030 -68.630 80.170 -68.620 ;
        RECT 79.950 -68.950 80.270 -68.630 ;
        RECT 73.070 -71.080 73.330 -70.760 ;
        RECT 73.130 -72.270 73.270 -71.080 ;
        RECT 73.130 -72.590 73.390 -72.270 ;
        RECT 73.130 -73.660 73.270 -72.590 ;
        RECT 73.040 -73.980 73.360 -73.660 ;
        RECT 80.030 -75.800 80.170 -68.950 ;
        RECT 79.950 -76.120 80.270 -75.800 ;
        RECT 82.700 -83.510 82.840 -61.230 ;
        RECT 91.880 -66.040 92.020 -48.780 ;
        RECT 94.540 -56.180 94.680 -33.900 ;
        RECT 102.150 -41.320 102.320 -27.260 ;
        RECT 106.300 -31.050 106.600 -30.650 ;
        RECT 106.380 -33.580 106.520 -31.050 ;
        RECT 106.290 -33.900 106.610 -33.580 ;
        RECT 102.110 -41.640 102.370 -41.320 ;
        RECT 96.790 -43.750 97.050 -43.430 ;
        RECT 96.850 -44.930 96.990 -43.750 ;
        RECT 103.640 -44.240 103.960 -43.920 ;
        RECT 96.810 -45.250 97.090 -44.930 ;
        RECT 96.850 -46.360 96.990 -45.250 ;
        RECT 96.760 -46.620 97.080 -46.360 ;
        RECT 103.720 -48.460 103.860 -44.240 ;
        RECT 103.630 -48.780 103.950 -48.460 ;
        RECT 94.450 -56.500 94.770 -56.180 ;
        RECT 94.540 -60.910 94.680 -56.500 ;
        RECT 94.450 -61.230 94.770 -60.910 ;
        RECT 91.800 -66.360 92.120 -66.040 ;
        RECT 91.870 -68.630 92.010 -68.620 ;
        RECT 91.790 -68.950 92.110 -68.630 ;
        RECT 84.890 -71.080 85.150 -70.760 ;
        RECT 84.950 -72.270 85.090 -71.080 ;
        RECT 84.950 -72.590 85.210 -72.270 ;
        RECT 84.950 -73.660 85.090 -72.590 ;
        RECT 84.860 -73.980 85.180 -73.660 ;
        RECT 91.870 -75.800 92.010 -68.950 ;
        RECT 91.790 -76.120 92.110 -75.800 ;
        RECT 94.540 -83.510 94.680 -61.230 ;
        RECT 103.720 -66.040 103.860 -48.780 ;
        RECT 106.380 -56.180 106.520 -33.900 ;
        RECT 114.280 -41.310 114.450 -26.630 ;
        RECT 118.170 -31.010 118.470 -30.610 ;
        RECT 118.250 -33.580 118.390 -31.010 ;
        RECT 118.160 -33.900 118.480 -33.580 ;
        RECT 114.240 -41.630 114.500 -41.310 ;
        RECT 108.630 -43.750 108.890 -43.430 ;
        RECT 108.690 -44.930 108.830 -43.750 ;
        RECT 115.510 -44.240 115.830 -43.920 ;
        RECT 108.650 -45.250 108.930 -44.930 ;
        RECT 108.690 -46.360 108.830 -45.250 ;
        RECT 108.600 -46.620 108.920 -46.360 ;
        RECT 115.590 -48.460 115.730 -44.240 ;
        RECT 115.500 -48.780 115.820 -48.460 ;
        RECT 106.290 -56.500 106.610 -56.180 ;
        RECT 106.380 -60.910 106.520 -56.500 ;
        RECT 106.290 -61.230 106.610 -60.910 ;
        RECT 103.640 -66.360 103.960 -66.040 ;
        RECT 103.710 -68.630 103.850 -68.620 ;
        RECT 103.630 -68.950 103.950 -68.630 ;
        RECT 96.730 -71.080 96.990 -70.760 ;
        RECT 96.790 -72.270 96.930 -71.080 ;
        RECT 96.790 -72.590 97.050 -72.270 ;
        RECT 96.790 -73.660 96.930 -72.590 ;
        RECT 96.700 -73.980 97.020 -73.660 ;
        RECT 103.710 -75.800 103.850 -68.950 ;
        RECT 103.630 -76.120 103.950 -75.800 ;
        RECT 106.380 -83.510 106.520 -61.230 ;
        RECT 115.590 -66.040 115.730 -48.780 ;
        RECT 118.250 -56.180 118.390 -33.900 ;
        RECT 125.910 -41.320 126.080 -26.130 ;
        RECT 130.040 -31.030 130.340 -30.630 ;
        RECT 130.120 -33.580 130.260 -31.030 ;
        RECT 130.030 -33.900 130.350 -33.580 ;
        RECT 125.870 -41.640 126.130 -41.320 ;
        RECT 120.500 -43.750 120.760 -43.430 ;
        RECT 120.560 -44.930 120.700 -43.750 ;
        RECT 127.380 -44.240 127.700 -43.920 ;
        RECT 120.520 -45.250 120.800 -44.930 ;
        RECT 120.560 -46.360 120.700 -45.250 ;
        RECT 120.470 -46.620 120.790 -46.360 ;
        RECT 127.460 -48.460 127.600 -44.240 ;
        RECT 127.370 -48.780 127.690 -48.460 ;
        RECT 118.160 -56.500 118.480 -56.180 ;
        RECT 118.250 -60.910 118.390 -56.500 ;
        RECT 118.160 -61.230 118.480 -60.910 ;
        RECT 115.510 -66.360 115.830 -66.040 ;
        RECT 115.580 -68.630 115.720 -68.620 ;
        RECT 115.500 -68.950 115.820 -68.630 ;
        RECT 108.570 -71.080 108.830 -70.760 ;
        RECT 108.630 -72.270 108.770 -71.080 ;
        RECT 108.630 -72.590 108.890 -72.270 ;
        RECT 108.630 -73.660 108.770 -72.590 ;
        RECT 108.540 -73.980 108.860 -73.660 ;
        RECT 115.580 -75.800 115.720 -68.950 ;
        RECT 115.500 -76.120 115.820 -75.800 ;
        RECT 118.250 -83.510 118.390 -61.230 ;
        RECT 127.460 -66.040 127.600 -48.780 ;
        RECT 130.120 -56.180 130.260 -33.900 ;
        RECT 135.370 -41.340 135.540 -25.660 ;
        RECT 139.050 -31.050 139.350 -30.650 ;
        RECT 139.130 -33.580 139.270 -31.050 ;
        RECT 139.040 -33.900 139.360 -33.580 ;
        RECT 135.300 -41.600 135.620 -41.340 ;
        RECT 132.370 -43.750 132.630 -43.430 ;
        RECT 132.430 -44.930 132.570 -43.750 ;
        RECT 136.390 -44.240 136.710 -43.920 ;
        RECT 132.390 -45.250 132.670 -44.930 ;
        RECT 132.430 -46.360 132.570 -45.250 ;
        RECT 132.340 -46.620 132.660 -46.360 ;
        RECT 136.470 -48.460 136.610 -44.240 ;
        RECT 136.380 -48.780 136.700 -48.460 ;
        RECT 130.030 -56.500 130.350 -56.180 ;
        RECT 130.120 -60.910 130.260 -56.500 ;
        RECT 130.030 -61.230 130.350 -60.910 ;
        RECT 127.380 -66.360 127.700 -66.040 ;
        RECT 127.450 -68.630 127.590 -68.620 ;
        RECT 127.370 -68.950 127.690 -68.630 ;
        RECT 120.440 -71.080 120.700 -70.760 ;
        RECT 120.500 -72.270 120.640 -71.080 ;
        RECT 120.500 -72.590 120.760 -72.270 ;
        RECT 120.500 -73.660 120.640 -72.590 ;
        RECT 120.410 -73.980 120.730 -73.660 ;
        RECT 127.450 -75.800 127.590 -68.950 ;
        RECT 127.370 -76.120 127.690 -75.800 ;
        RECT 130.120 -83.510 130.260 -61.230 ;
        RECT 136.470 -66.040 136.610 -48.780 ;
        RECT 139.130 -56.180 139.270 -33.900 ;
        RECT 141.380 -43.750 141.640 -43.430 ;
        RECT 141.440 -44.930 141.580 -43.750 ;
        RECT 141.400 -45.250 141.680 -44.930 ;
        RECT 141.440 -46.360 141.580 -45.250 ;
        RECT 141.350 -46.620 141.670 -46.360 ;
        RECT 139.040 -56.500 139.360 -56.180 ;
        RECT 139.130 -60.910 139.270 -56.500 ;
        RECT 139.040 -61.230 139.360 -60.910 ;
        RECT 136.390 -66.360 136.710 -66.040 ;
        RECT 136.460 -68.630 136.600 -68.620 ;
        RECT 136.380 -68.950 136.700 -68.630 ;
        RECT 132.310 -71.080 132.570 -70.760 ;
        RECT 132.370 -72.270 132.510 -71.080 ;
        RECT 132.370 -72.590 132.630 -72.270 ;
        RECT 132.370 -73.660 132.510 -72.590 ;
        RECT 132.280 -73.980 132.600 -73.660 ;
        RECT 136.460 -75.800 136.600 -68.950 ;
        RECT 136.380 -76.120 136.700 -75.800 ;
        RECT 139.130 -83.510 139.270 -61.230 ;
        RECT 141.320 -71.080 141.580 -70.760 ;
        RECT 141.380 -72.270 141.520 -71.080 ;
        RECT 141.380 -72.590 141.640 -72.270 ;
        RECT 141.380 -73.660 141.520 -72.590 ;
        RECT 141.290 -73.980 141.610 -73.660 ;
        RECT -35.250 -83.830 -34.930 -83.510 ;
        RECT -23.750 -83.830 -23.430 -83.510 ;
        RECT -11.930 -83.830 -11.610 -83.510 ;
        RECT -0.120 -83.830 0.200 -83.510 ;
        RECT 11.690 -83.830 12.010 -83.510 ;
        RECT 23.510 -83.830 23.830 -83.510 ;
        RECT 35.330 -83.830 35.650 -83.510 ;
        RECT 47.150 -83.830 47.470 -83.510 ;
        RECT 58.970 -83.830 59.290 -83.510 ;
        RECT 70.790 -83.830 71.110 -83.510 ;
        RECT 82.610 -83.830 82.930 -83.510 ;
        RECT 94.450 -83.830 94.770 -83.510 ;
        RECT 106.290 -83.830 106.610 -83.510 ;
        RECT 118.160 -83.830 118.480 -83.510 ;
        RECT 130.030 -83.830 130.350 -83.510 ;
        RECT 139.040 -83.830 139.360 -83.510 ;
        RECT -35.160 -86.240 -35.020 -83.830 ;
        RECT -23.660 -86.240 -23.520 -83.830 ;
        RECT -11.840 -86.240 -11.700 -83.830 ;
        RECT -0.030 -86.240 0.110 -83.830 ;
        RECT 11.780 -86.240 11.920 -83.830 ;
        RECT 23.600 -86.240 23.740 -83.830 ;
        RECT 35.420 -86.240 35.560 -83.830 ;
        RECT 47.240 -86.240 47.380 -83.830 ;
        RECT 59.060 -86.240 59.200 -83.830 ;
        RECT 70.880 -86.240 71.020 -83.830 ;
        RECT 82.700 -86.240 82.840 -83.830 ;
        RECT 94.540 -86.240 94.680 -83.830 ;
        RECT 106.380 -86.240 106.520 -83.830 ;
        RECT 118.250 -86.240 118.390 -83.830 ;
        RECT 130.120 -86.240 130.260 -83.830 ;
        RECT 139.130 -86.240 139.270 -83.830 ;
      LAYER via2 ;
        RECT -43.140 50.310 -42.840 50.610 ;
        RECT 5.240 50.390 5.540 50.690 ;
        RECT 11.000 50.390 11.300 50.690 ;
        RECT 16.750 50.390 17.050 50.690 ;
        RECT 22.480 50.390 22.780 50.690 ;
        RECT 28.240 50.390 28.540 50.690 ;
        RECT 33.980 50.390 34.280 50.690 ;
        RECT 39.730 50.390 40.030 50.690 ;
        RECT 45.480 50.390 45.780 50.690 ;
        RECT 51.230 50.390 51.530 50.690 ;
        RECT 56.990 50.390 57.290 50.690 ;
        RECT 62.740 50.380 63.040 50.680 ;
        RECT 68.480 50.390 68.780 50.690 ;
        RECT 74.230 50.390 74.530 50.690 ;
        RECT 79.980 50.390 80.280 50.690 ;
        RECT 85.720 50.390 86.020 50.690 ;
        RECT 91.470 50.390 91.770 50.690 ;
        RECT 5.960 -6.370 6.260 -6.070 ;
        RECT -41.800 -20.640 -41.500 -20.340 ;
        RECT -0.350 -20.600 -0.050 -20.300 ;
        RECT -43.140 -30.930 -42.840 -30.630 ;
        RECT 11.710 -7.640 12.010 -7.340 ;
        RECT 17.510 -9.010 17.810 -8.710 ;
        RECT 8.110 -23.500 8.410 -23.200 ;
        RECT 23.210 -10.180 23.510 -9.880 ;
        RECT 19.600 -23.510 19.900 -23.210 ;
        RECT 28.960 -11.430 29.260 -11.130 ;
        RECT 34.710 -12.880 35.010 -12.580 ;
        RECT 31.030 -23.520 31.330 -23.220 ;
        RECT 40.450 -14.100 40.750 -13.800 ;
        RECT 46.210 -14.980 46.510 -14.680 ;
        RECT 42.600 -23.530 42.900 -23.230 ;
        RECT 51.960 -15.810 52.260 -15.510 ;
        RECT 57.710 -16.590 58.010 -16.290 ;
        RECT 54.000 -23.510 54.300 -23.210 ;
        RECT 63.460 -17.450 63.760 -17.150 ;
        RECT 69.210 -18.250 69.510 -17.950 ;
        RECT 65.680 -23.510 65.980 -23.210 ;
        RECT 74.960 -19.050 75.260 -18.750 ;
        RECT 80.710 -19.700 81.010 -19.400 ;
        RECT 77.130 -23.510 77.430 -23.210 ;
        RECT 86.460 -20.840 86.760 -20.540 ;
        RECT 92.210 -21.730 92.510 -21.430 ;
        RECT 88.700 -23.490 89.000 -23.190 ;
        RECT 7.350 -24.490 7.650 -24.190 ;
        RECT 8.900 -24.490 9.200 -24.190 ;
        RECT 18.850 -24.490 19.150 -24.190 ;
        RECT 20.400 -24.490 20.700 -24.190 ;
        RECT 30.350 -24.490 30.650 -24.190 ;
        RECT 31.890 -24.490 32.190 -24.190 ;
        RECT 41.820 -24.490 42.120 -24.190 ;
        RECT 43.410 -24.500 43.710 -24.200 ;
        RECT 53.340 -24.490 53.640 -24.190 ;
        RECT 54.890 -24.490 55.190 -24.190 ;
        RECT 64.850 -24.500 65.150 -24.200 ;
        RECT 66.380 -24.500 66.680 -24.200 ;
        RECT 76.360 -24.490 76.660 -24.190 ;
        RECT 77.890 -24.490 78.190 -24.190 ;
        RECT 87.850 -24.480 88.150 -24.180 ;
        RECT 89.370 -24.490 89.670 -24.190 ;
        RECT 4.660 -25.260 4.960 -24.960 ;
        RECT 11.590 -25.190 11.890 -24.890 ;
        RECT 16.150 -25.180 16.450 -24.880 ;
        RECT 23.080 -25.230 23.380 -24.930 ;
        RECT 27.670 -25.240 27.970 -24.940 ;
        RECT 34.590 -25.220 34.890 -24.920 ;
        RECT 39.170 -25.240 39.470 -24.940 ;
        RECT 46.080 -25.260 46.380 -24.960 ;
        RECT 50.660 -25.200 50.960 -24.900 ;
        RECT 57.590 -25.220 57.890 -24.920 ;
        RECT 62.160 -25.180 62.460 -24.880 ;
        RECT 69.080 -25.220 69.380 -24.920 ;
        RECT 73.660 -25.220 73.960 -24.920 ;
        RECT 80.580 -25.250 80.880 -24.950 ;
        RECT 85.160 -25.230 85.460 -24.930 ;
        RECT 92.070 -25.200 92.350 -24.920 ;
        RECT -35.240 -30.970 -34.940 -30.670 ;
        RECT -23.740 -30.970 -23.440 -30.670 ;
        RECT -0.110 -31.010 0.190 -30.710 ;
        RECT 11.700 -30.990 12.000 -30.690 ;
        RECT 23.520 -31.000 23.820 -30.700 ;
        RECT 35.340 -31.000 35.640 -30.700 ;
        RECT 47.160 -30.970 47.460 -30.670 ;
        RECT 58.980 -31.000 59.280 -30.700 ;
        RECT 70.800 -31.000 71.100 -30.700 ;
        RECT 82.620 -30.980 82.920 -30.680 ;
        RECT 94.460 -30.990 94.760 -30.690 ;
        RECT 106.300 -31.000 106.600 -30.700 ;
        RECT 118.170 -30.960 118.470 -30.660 ;
        RECT 130.040 -30.980 130.340 -30.680 ;
        RECT 139.050 -31.000 139.350 -30.700 ;
  END
END Integrated_bitcell_with_dummy_cells
END LIBRARY

