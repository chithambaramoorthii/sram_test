magic
tech sky130B
timestamp 1662734547
<< nwell >>
rect 225 5055 304 5059
rect 321 5055 395 5059
rect 412 5055 660 5059
rect 690 5055 755 5059
rect 785 5055 873 5059
rect 903 5055 965 5059
rect 995 5055 1235 5059
rect 1265 5055 1328 5059
rect 1358 5055 1449 5059
rect 1479 5055 1543 5059
rect 1573 5055 1810 5059
rect 1840 5055 1907 5059
rect 1937 5055 2024 5059
rect 2054 5055 2116 5059
rect 2146 5055 2376 5059
rect 2734 5055 2959 5059
rect 3317 5055 3526 5059
rect 3884 5055 4103 5059
rect 4461 5055 4674 5059
rect 5032 5055 5258 5059
rect 5616 5055 5838 5059
rect 6196 5055 6413 5059
rect 6771 5055 6989 5059
rect 7347 5055 7563 5059
rect 7921 5055 8137 5059
rect 8495 5055 8714 5059
rect 9072 5055 9287 5059
rect 1095 5034 1135 5055
rect 1670 5034 1710 5055
rect 2243 5034 2283 5055
rect 2819 5034 2859 5055
rect 3393 5034 3433 5055
rect 3968 5034 4008 5055
rect 4543 5034 4583 5055
rect 5118 5034 5158 5055
rect 5694 5034 5734 5055
rect 6269 5033 6309 5055
rect 6843 5034 6883 5055
rect 7418 5034 7458 5055
rect 7993 5034 8033 5055
rect 8567 5034 8607 5055
rect 9142 5034 9182 5055
rect 604 -1408 609 -1395
rect 601 -1412 618 -1408
rect 797 -2200 827 -2183
rect 1340 -2210 1416 -2174
rect 1915 -2210 1991 -2174
rect 2490 -2210 2566 -2174
rect 3065 -2210 3141 -2174
rect 3640 -2210 3716 -2174
rect 4215 -2210 4291 -2174
rect 4790 -2210 4866 -2174
rect 5365 -2210 5441 -2174
rect 5940 -2210 6016 -2174
rect 6515 -2210 6591 -2174
rect 7090 -2210 7166 -2174
rect 7665 -2210 7741 -2174
rect 8240 -2210 8316 -2174
rect 8815 -2184 8891 -2174
rect 8904 -2184 8940 -2183
rect 8815 -2200 8940 -2184
rect 8815 -2201 8935 -2200
rect 8815 -2210 8891 -2201
rect 585 -2256 589 -2255
rect 225 -2454 589 -2256
rect 1064 -2454 1739 -2256
rect 2214 -2454 2889 -2256
rect 3364 -2454 4039 -2256
rect 4514 -2454 5189 -2256
rect 5664 -2454 6339 -2256
rect 6814 -2454 7489 -2256
rect 7964 -2454 8639 -2256
rect 9114 -2454 9466 -2256
rect -3516 -3121 -3502 -3117
<< pwell >>
rect 225 4109 470 4482
rect 225 3583 231 3597
rect 224 3342 230 3356
rect 225 3101 231 3115
rect 224 2860 230 2874
rect 225 2579 231 2593
rect 225 2338 231 2352
rect 225 2097 231 2111
rect 225 1856 231 1870
rect 225 1615 231 1629
rect 225 1374 231 1388
rect 225 1133 231 1147
rect 225 892 231 906
rect 225 610 231 624
rect 225 369 231 383
rect 225 128 231 142
rect 225 -1866 228 -1852
rect 225 -1913 228 -1899
rect 812 -1913 829 -1896
rect 1375 -1924 1416 -1888
rect 1950 -1924 1991 -1888
rect 2525 -1924 2566 -1888
rect 3100 -1924 3141 -1888
rect 3675 -1924 3716 -1888
rect 4250 -1924 4291 -1888
rect 4825 -1924 4866 -1888
rect 5400 -1924 5441 -1888
rect 5975 -1924 6016 -1888
rect 6550 -1924 6591 -1888
rect 7125 -1924 7166 -1888
rect 7700 -1924 7741 -1888
rect 8275 -1924 8316 -1888
rect 8850 -1924 8891 -1888
rect 9411 -1924 9452 -1888
rect 225 -1964 228 -1950
rect 225 -2052 228 -2038
rect 589 -2454 1064 -2256
rect 1739 -2454 2214 -2256
rect 2889 -2454 3364 -2256
rect 4039 -2454 4514 -2256
rect 5189 -2454 5664 -2256
rect 6339 -2454 6814 -2256
rect 7489 -2454 7964 -2256
rect 8639 -2454 9114 -2256
rect 14196 -4434 14214 -4417
rect -889 -4562 -860 -4539
rect 14179 -4589 14214 -4572
rect 14196 -7169 14214 -7152
rect 14196 -7321 14214 -7304
<< nmos >>
rect 646 -2387 710 -2372
rect 943 -2387 1007 -2372
rect 1796 -2392 1860 -2377
rect 2093 -2392 2157 -2377
rect 2946 -2392 3010 -2377
rect 3243 -2392 3307 -2377
rect 4096 -2392 4160 -2377
rect 4393 -2392 4457 -2377
rect 5246 -2392 5310 -2377
rect 5543 -2392 5607 -2377
rect 6396 -2392 6460 -2377
rect 6693 -2392 6757 -2377
rect 7546 -2392 7610 -2377
rect 7843 -2392 7907 -2377
rect 8696 -2392 8760 -2377
rect 8993 -2392 9057 -2377
<< pmos >>
rect 518 -2387 560 -2372
rect 1093 -2387 1135 -2372
rect 1668 -2392 1710 -2377
rect 2243 -2392 2285 -2377
rect 2818 -2392 2860 -2377
rect 3393 -2392 3435 -2377
rect 3968 -2392 4010 -2377
rect 4543 -2392 4585 -2377
rect 5118 -2392 5160 -2377
rect 5693 -2392 5735 -2377
rect 6268 -2392 6310 -2377
rect 6843 -2392 6885 -2377
rect 7418 -2392 7460 -2377
rect 7993 -2392 8035 -2377
rect 8568 -2392 8610 -2377
rect 9143 -2392 9185 -2377
<< ndiff >>
rect 646 -2348 710 -2342
rect 646 -2365 668 -2348
rect 685 -2365 710 -2348
rect 943 -2347 1007 -2342
rect 646 -2372 710 -2365
rect 646 -2395 710 -2387
rect 646 -2412 669 -2395
rect 686 -2412 710 -2395
rect 943 -2364 967 -2347
rect 984 -2364 1007 -2347
rect 943 -2372 1007 -2364
rect 943 -2394 1007 -2387
rect 646 -2417 710 -2412
rect 943 -2411 968 -2394
rect 985 -2411 1007 -2394
rect 943 -2417 1007 -2411
rect 1796 -2352 1860 -2347
rect 1796 -2369 1819 -2352
rect 1836 -2369 1860 -2352
rect 2093 -2352 2157 -2347
rect 1796 -2377 1860 -2369
rect 1796 -2400 1860 -2392
rect 1796 -2417 1818 -2400
rect 1835 -2417 1860 -2400
rect 2093 -2369 2117 -2352
rect 2134 -2369 2157 -2352
rect 2093 -2377 2157 -2369
rect 2093 -2400 2157 -2392
rect 1796 -2422 1860 -2417
rect 2093 -2417 2118 -2400
rect 2135 -2417 2157 -2400
rect 2093 -2422 2157 -2417
rect 2946 -2352 3010 -2347
rect 2946 -2369 2969 -2352
rect 2986 -2369 3010 -2352
rect 3243 -2352 3307 -2347
rect 2946 -2377 3010 -2369
rect 2946 -2400 3010 -2392
rect 2946 -2417 2968 -2400
rect 2985 -2417 3010 -2400
rect 3243 -2369 3267 -2352
rect 3284 -2369 3307 -2352
rect 3243 -2377 3307 -2369
rect 3243 -2400 3307 -2392
rect 2946 -2422 3010 -2417
rect 3243 -2418 3268 -2400
rect 3285 -2418 3307 -2400
rect 3243 -2422 3307 -2418
rect 4096 -2352 4160 -2347
rect 4096 -2369 4119 -2352
rect 4136 -2369 4160 -2352
rect 4393 -2352 4457 -2347
rect 4096 -2377 4160 -2369
rect 4096 -2400 4160 -2392
rect 4096 -2417 4118 -2400
rect 4135 -2417 4160 -2400
rect 4393 -2369 4417 -2352
rect 4434 -2369 4457 -2352
rect 4393 -2377 4457 -2369
rect 4393 -2400 4457 -2392
rect 4096 -2422 4160 -2417
rect 4393 -2417 4418 -2400
rect 4435 -2417 4457 -2400
rect 4393 -2422 4457 -2417
rect 5246 -2352 5310 -2347
rect 5246 -2369 5269 -2352
rect 5286 -2369 5310 -2352
rect 5543 -2352 5607 -2347
rect 5246 -2377 5310 -2369
rect 5246 -2400 5310 -2392
rect 5246 -2417 5268 -2400
rect 5285 -2417 5310 -2400
rect 5543 -2369 5567 -2352
rect 5584 -2369 5607 -2352
rect 5543 -2377 5607 -2369
rect 5543 -2400 5607 -2392
rect 5246 -2422 5310 -2417
rect 5543 -2417 5568 -2400
rect 5585 -2417 5607 -2400
rect 5543 -2422 5607 -2417
rect 6396 -2352 6460 -2347
rect 6396 -2369 6419 -2352
rect 6436 -2369 6460 -2352
rect 6693 -2352 6757 -2347
rect 6396 -2377 6460 -2369
rect 6396 -2400 6460 -2392
rect 6396 -2417 6418 -2400
rect 6435 -2417 6460 -2400
rect 6693 -2369 6717 -2352
rect 6734 -2369 6757 -2352
rect 6693 -2377 6757 -2369
rect 6693 -2400 6757 -2392
rect 6396 -2422 6460 -2417
rect 6693 -2417 6718 -2400
rect 6735 -2417 6757 -2400
rect 6693 -2422 6757 -2417
rect 7546 -2352 7610 -2347
rect 7546 -2369 7569 -2352
rect 7586 -2369 7610 -2352
rect 7843 -2352 7907 -2347
rect 7546 -2377 7610 -2369
rect 7546 -2400 7610 -2392
rect 7546 -2417 7568 -2400
rect 7585 -2417 7610 -2400
rect 7843 -2369 7867 -2352
rect 7884 -2369 7907 -2352
rect 7843 -2377 7907 -2369
rect 7843 -2400 7907 -2392
rect 7546 -2422 7610 -2417
rect 7843 -2417 7868 -2400
rect 7885 -2417 7907 -2400
rect 7843 -2422 7907 -2417
rect 8696 -2352 8760 -2347
rect 8696 -2369 8719 -2352
rect 8736 -2369 8760 -2352
rect 8993 -2352 9057 -2347
rect 8696 -2377 8760 -2369
rect 8696 -2400 8760 -2392
rect 8696 -2417 8718 -2400
rect 8735 -2417 8760 -2400
rect 8993 -2369 9017 -2352
rect 9034 -2369 9057 -2352
rect 8993 -2377 9057 -2369
rect 8993 -2400 9057 -2392
rect 8696 -2422 8760 -2417
rect 8993 -2417 9018 -2400
rect 9035 -2417 9057 -2400
rect 8993 -2422 9057 -2417
<< pdiff >>
rect 518 -2347 560 -2338
rect 518 -2364 531 -2347
rect 548 -2364 560 -2347
rect 518 -2372 560 -2364
rect 518 -2395 560 -2387
rect 518 -2412 531 -2395
rect 548 -2412 560 -2395
rect 518 -2417 560 -2412
rect 1093 -2347 1135 -2342
rect 1093 -2364 1105 -2347
rect 1122 -2364 1135 -2347
rect 1668 -2352 1710 -2347
rect 1093 -2372 1135 -2364
rect 1093 -2394 1135 -2387
rect 1093 -2411 1105 -2394
rect 1122 -2411 1135 -2394
rect 1668 -2369 1681 -2352
rect 1698 -2369 1710 -2352
rect 1668 -2377 1710 -2369
rect 1668 -2400 1710 -2392
rect 1093 -2421 1135 -2411
rect 1668 -2417 1681 -2400
rect 1698 -2417 1710 -2400
rect 1668 -2426 1710 -2417
rect 2243 -2352 2285 -2347
rect 2243 -2369 2255 -2352
rect 2272 -2369 2285 -2352
rect 2818 -2352 2860 -2347
rect 2243 -2377 2285 -2369
rect 2243 -2400 2285 -2392
rect 2818 -2369 2831 -2352
rect 2848 -2369 2860 -2352
rect 2818 -2377 2860 -2369
rect 2818 -2400 2860 -2392
rect 2243 -2417 2255 -2400
rect 2272 -2417 2285 -2400
rect 2243 -2426 2285 -2417
rect 2818 -2417 2831 -2400
rect 2848 -2417 2860 -2400
rect 2818 -2426 2860 -2417
rect 3393 -2352 3435 -2347
rect 3393 -2369 3405 -2352
rect 3422 -2369 3435 -2352
rect 3968 -2352 4010 -2347
rect 3393 -2377 3435 -2369
rect 3393 -2400 3435 -2392
rect 3968 -2369 3981 -2352
rect 3998 -2369 4010 -2352
rect 3968 -2377 4010 -2369
rect 3968 -2400 4010 -2392
rect 3393 -2417 3405 -2400
rect 3422 -2417 3435 -2400
rect 3393 -2426 3435 -2417
rect 3968 -2417 3981 -2400
rect 3998 -2417 4010 -2400
rect 3968 -2426 4010 -2417
rect 4543 -2352 4585 -2347
rect 4543 -2369 4555 -2352
rect 4572 -2369 4585 -2352
rect 5118 -2352 5160 -2347
rect 4543 -2377 4585 -2369
rect 4543 -2400 4585 -2392
rect 5118 -2369 5131 -2352
rect 5148 -2369 5160 -2352
rect 5118 -2377 5160 -2369
rect 5118 -2400 5160 -2392
rect 4543 -2417 4555 -2400
rect 4572 -2417 4585 -2400
rect 4543 -2426 4585 -2417
rect 5118 -2417 5131 -2400
rect 5148 -2417 5160 -2400
rect 5118 -2426 5160 -2417
rect 5693 -2352 5735 -2347
rect 5693 -2369 5705 -2352
rect 5722 -2369 5735 -2352
rect 6268 -2352 6310 -2347
rect 5693 -2377 5735 -2369
rect 5693 -2400 5735 -2392
rect 6268 -2369 6281 -2352
rect 6298 -2369 6310 -2352
rect 6268 -2377 6310 -2369
rect 6268 -2400 6310 -2392
rect 5693 -2417 5705 -2400
rect 5722 -2417 5735 -2400
rect 5693 -2426 5735 -2417
rect 6268 -2417 6281 -2400
rect 6298 -2417 6310 -2400
rect 6268 -2426 6310 -2417
rect 6843 -2352 6885 -2347
rect 6843 -2369 6855 -2352
rect 6872 -2369 6885 -2352
rect 7418 -2352 7460 -2347
rect 6843 -2377 6885 -2369
rect 6843 -2400 6885 -2392
rect 7418 -2369 7431 -2352
rect 7448 -2369 7460 -2352
rect 7418 -2377 7460 -2369
rect 7418 -2400 7460 -2392
rect 6843 -2417 6855 -2400
rect 6872 -2417 6885 -2400
rect 6843 -2426 6885 -2417
rect 7418 -2417 7431 -2400
rect 7448 -2417 7460 -2400
rect 7418 -2426 7460 -2417
rect 7993 -2352 8035 -2347
rect 7993 -2369 8005 -2352
rect 8022 -2369 8035 -2352
rect 8568 -2352 8610 -2347
rect 7993 -2377 8035 -2369
rect 7993 -2400 8035 -2392
rect 8568 -2369 8581 -2352
rect 8598 -2369 8610 -2352
rect 8568 -2377 8610 -2369
rect 8568 -2400 8610 -2392
rect 7993 -2417 8005 -2400
rect 8022 -2417 8035 -2400
rect 7993 -2426 8035 -2417
rect 8568 -2417 8581 -2400
rect 8598 -2417 8610 -2400
rect 8568 -2426 8610 -2417
rect 9143 -2352 9185 -2347
rect 9143 -2369 9155 -2352
rect 9172 -2369 9185 -2352
rect 9143 -2377 9185 -2369
rect 9143 -2400 9185 -2392
rect 9143 -2417 9155 -2400
rect 9172 -2417 9185 -2400
rect 9143 -2426 9185 -2417
<< ndiffc >>
rect 668 -2365 685 -2348
rect 669 -2412 686 -2395
rect 967 -2364 984 -2347
rect 968 -2411 985 -2394
rect 1819 -2369 1836 -2352
rect 1818 -2417 1835 -2400
rect 2117 -2369 2134 -2352
rect 2118 -2417 2135 -2400
rect 2969 -2369 2986 -2352
rect 2968 -2417 2985 -2400
rect 3267 -2369 3284 -2352
rect 3268 -2418 3285 -2400
rect 4119 -2369 4136 -2352
rect 4118 -2417 4135 -2400
rect 4417 -2369 4434 -2352
rect 4418 -2417 4435 -2400
rect 5269 -2369 5286 -2352
rect 5268 -2417 5285 -2400
rect 5567 -2369 5584 -2352
rect 5568 -2417 5585 -2400
rect 6419 -2369 6436 -2352
rect 6418 -2417 6435 -2400
rect 6717 -2369 6734 -2352
rect 6718 -2417 6735 -2400
rect 7569 -2369 7586 -2352
rect 7568 -2417 7585 -2400
rect 7867 -2369 7884 -2352
rect 7868 -2417 7885 -2400
rect 8719 -2369 8736 -2352
rect 8718 -2417 8735 -2400
rect 9017 -2369 9034 -2352
rect 9018 -2417 9035 -2400
<< pdiffc >>
rect 531 -2364 548 -2347
rect 531 -2412 548 -2395
rect 1105 -2364 1122 -2347
rect 1105 -2411 1122 -2394
rect 1681 -2369 1698 -2352
rect 1681 -2417 1698 -2400
rect 2255 -2369 2272 -2352
rect 2831 -2369 2848 -2352
rect 2255 -2417 2272 -2400
rect 2831 -2417 2848 -2400
rect 3405 -2369 3422 -2352
rect 3981 -2369 3998 -2352
rect 3405 -2417 3422 -2400
rect 3981 -2417 3998 -2400
rect 4555 -2369 4572 -2352
rect 5131 -2369 5148 -2352
rect 4555 -2417 4572 -2400
rect 5131 -2417 5148 -2400
rect 5705 -2369 5722 -2352
rect 6281 -2369 6298 -2352
rect 5705 -2417 5722 -2400
rect 6281 -2417 6298 -2400
rect 6855 -2369 6872 -2352
rect 7431 -2369 7448 -2352
rect 6855 -2417 6872 -2400
rect 7431 -2417 7448 -2400
rect 8005 -2369 8022 -2352
rect 8581 -2369 8598 -2352
rect 8005 -2417 8022 -2400
rect 8581 -2417 8598 -2400
rect 9155 -2369 9172 -2352
rect 9155 -2417 9172 -2400
<< psubdiff >>
rect 800 -1896 841 -1888
rect 800 -1913 812 -1896
rect 829 -1913 841 -1896
rect 800 -1924 841 -1913
rect 1375 -1896 1416 -1888
rect 1375 -1913 1387 -1896
rect 1404 -1913 1416 -1896
rect 1375 -1924 1416 -1913
rect 1950 -1896 1991 -1888
rect 1950 -1913 1962 -1896
rect 1979 -1913 1991 -1896
rect 1950 -1924 1991 -1913
rect 2525 -1896 2566 -1888
rect 2525 -1913 2537 -1896
rect 2554 -1913 2566 -1896
rect 2525 -1924 2566 -1913
rect 3100 -1896 3141 -1888
rect 3100 -1913 3112 -1896
rect 3129 -1913 3141 -1896
rect 3100 -1924 3141 -1913
rect 3675 -1896 3716 -1888
rect 3675 -1913 3687 -1896
rect 3704 -1913 3716 -1896
rect 3675 -1924 3716 -1913
rect 4250 -1896 4291 -1888
rect 4250 -1913 4262 -1896
rect 4279 -1913 4291 -1896
rect 4250 -1924 4291 -1913
rect 4825 -1896 4866 -1888
rect 4825 -1913 4837 -1896
rect 4854 -1913 4866 -1896
rect 4825 -1924 4866 -1913
rect 5400 -1896 5441 -1888
rect 5400 -1913 5412 -1896
rect 5429 -1913 5441 -1896
rect 5400 -1924 5441 -1913
rect 5975 -1896 6016 -1888
rect 5975 -1913 5987 -1896
rect 6004 -1913 6016 -1896
rect 5975 -1924 6016 -1913
rect 6550 -1896 6591 -1888
rect 6550 -1913 6562 -1896
rect 6579 -1913 6591 -1896
rect 6550 -1924 6591 -1913
rect 7125 -1896 7166 -1888
rect 7125 -1913 7137 -1896
rect 7154 -1913 7166 -1896
rect 7125 -1924 7166 -1913
rect 7700 -1896 7741 -1888
rect 7700 -1913 7712 -1896
rect 7729 -1913 7741 -1896
rect 7700 -1924 7741 -1913
rect 8275 -1896 8316 -1888
rect 8275 -1913 8287 -1896
rect 8304 -1913 8316 -1896
rect 8275 -1924 8316 -1913
rect 8850 -1896 8891 -1888
rect 8850 -1913 8862 -1896
rect 8879 -1913 8891 -1896
rect 8850 -1924 8891 -1913
rect 9411 -1896 9452 -1888
rect 9411 -1913 9423 -1896
rect 9440 -1913 9452 -1896
rect 9411 -1924 9452 -1913
rect 805 -2326 846 -2318
rect 805 -2343 817 -2326
rect 834 -2343 846 -2326
rect 1954 -2327 1995 -2319
rect 805 -2354 846 -2343
rect 1954 -2344 1966 -2327
rect 1983 -2344 1995 -2327
rect 1954 -2355 1995 -2344
rect 3097 -2328 3138 -2320
rect 3097 -2345 3109 -2328
rect 3126 -2345 3138 -2328
rect 3097 -2356 3138 -2345
rect 4254 -2329 4295 -2321
rect 4254 -2346 4266 -2329
rect 4283 -2346 4295 -2329
rect 4254 -2357 4295 -2346
rect 5394 -2327 5435 -2319
rect 5394 -2344 5406 -2327
rect 5423 -2344 5435 -2327
rect 5394 -2355 5435 -2344
rect 6562 -2327 6603 -2319
rect 6562 -2344 6574 -2327
rect 6591 -2344 6603 -2327
rect 6562 -2355 6603 -2344
rect 7707 -2327 7748 -2319
rect 7707 -2344 7719 -2327
rect 7736 -2344 7748 -2327
rect 7707 -2355 7748 -2344
rect 8864 -2325 8905 -2317
rect 8864 -2342 8876 -2325
rect 8893 -2342 8905 -2325
rect 8864 -2353 8905 -2342
<< nsubdiff >>
rect 800 -2183 841 -2173
rect 800 -2200 812 -2183
rect 829 -2200 841 -2183
rect 800 -2209 841 -2200
rect 1375 -2184 1416 -2174
rect 1375 -2201 1387 -2184
rect 1404 -2201 1416 -2184
rect 1375 -2210 1416 -2201
rect 1950 -2184 1991 -2174
rect 1950 -2201 1962 -2184
rect 1979 -2201 1991 -2184
rect 1950 -2210 1991 -2201
rect 2525 -2184 2566 -2174
rect 2525 -2201 2537 -2184
rect 2554 -2201 2566 -2184
rect 2525 -2210 2566 -2201
rect 3100 -2184 3141 -2174
rect 3100 -2201 3112 -2184
rect 3129 -2201 3141 -2184
rect 3100 -2210 3141 -2201
rect 3675 -2184 3716 -2174
rect 3675 -2201 3687 -2184
rect 3704 -2201 3716 -2184
rect 3675 -2210 3716 -2201
rect 4250 -2184 4291 -2174
rect 4250 -2201 4262 -2184
rect 4279 -2201 4291 -2184
rect 4250 -2210 4291 -2201
rect 4825 -2184 4866 -2174
rect 4825 -2201 4837 -2184
rect 4854 -2201 4866 -2184
rect 4825 -2210 4866 -2201
rect 5400 -2184 5441 -2174
rect 5400 -2201 5412 -2184
rect 5429 -2201 5441 -2184
rect 5400 -2210 5441 -2201
rect 5975 -2184 6016 -2174
rect 5975 -2201 5987 -2184
rect 6004 -2201 6016 -2184
rect 5975 -2210 6016 -2201
rect 6550 -2184 6591 -2174
rect 6550 -2201 6562 -2184
rect 6579 -2201 6591 -2184
rect 6550 -2210 6591 -2201
rect 7125 -2184 7166 -2174
rect 7125 -2201 7137 -2184
rect 7154 -2201 7166 -2184
rect 7125 -2210 7166 -2201
rect 7700 -2184 7741 -2174
rect 7700 -2201 7712 -2184
rect 7729 -2201 7741 -2184
rect 7700 -2210 7741 -2201
rect 8275 -2184 8316 -2174
rect 8275 -2201 8287 -2184
rect 8304 -2201 8316 -2184
rect 8275 -2210 8316 -2201
rect 8850 -2184 8891 -2174
rect 8850 -2201 8862 -2184
rect 8879 -2201 8891 -2184
rect 8850 -2210 8891 -2201
<< psubdiffcont >>
rect 812 -1913 829 -1896
rect 1387 -1913 1404 -1896
rect 1962 -1913 1979 -1896
rect 2537 -1913 2554 -1896
rect 3112 -1913 3129 -1896
rect 3687 -1913 3704 -1896
rect 4262 -1913 4279 -1896
rect 4837 -1913 4854 -1896
rect 5412 -1913 5429 -1896
rect 5987 -1913 6004 -1896
rect 6562 -1913 6579 -1896
rect 7137 -1913 7154 -1896
rect 7712 -1913 7729 -1896
rect 8287 -1913 8304 -1896
rect 8862 -1913 8879 -1896
rect 9423 -1913 9440 -1896
rect 817 -2343 834 -2326
rect 1966 -2344 1983 -2327
rect 3109 -2345 3126 -2328
rect 4266 -2346 4283 -2329
rect 5406 -2344 5423 -2327
rect 6574 -2344 6591 -2327
rect 7719 -2344 7736 -2327
rect 8876 -2342 8893 -2325
<< nsubdiffcont >>
rect 812 -2200 829 -2183
rect 1387 -2201 1404 -2184
rect 1962 -2201 1979 -2184
rect 2537 -2201 2554 -2184
rect 3112 -2201 3129 -2184
rect 3687 -2201 3704 -2184
rect 4262 -2201 4279 -2184
rect 4837 -2201 4854 -2184
rect 5412 -2201 5429 -2184
rect 5987 -2201 6004 -2184
rect 6562 -2201 6579 -2184
rect 7137 -2201 7154 -2184
rect 7712 -2201 7729 -2184
rect 8287 -2201 8304 -2184
rect 8862 -2201 8879 -2184
<< poly >>
rect 464 -2372 497 -2364
rect 733 -2371 766 -2363
rect 733 -2372 741 -2371
rect 464 -2389 472 -2372
rect 489 -2387 518 -2372
rect 560 -2387 573 -2372
rect 633 -2387 646 -2372
rect 710 -2387 741 -2372
rect 489 -2389 497 -2387
rect 464 -2397 497 -2389
rect 733 -2388 741 -2387
rect 758 -2388 766 -2371
rect 733 -2396 766 -2388
rect 887 -2371 920 -2363
rect 887 -2388 895 -2371
rect 912 -2372 920 -2371
rect 1156 -2370 1189 -2362
rect 1156 -2372 1164 -2370
rect 912 -2387 943 -2372
rect 1007 -2387 1020 -2372
rect 1080 -2387 1093 -2372
rect 1135 -2387 1164 -2372
rect 1181 -2387 1189 -2370
rect 912 -2388 920 -2387
rect 887 -2396 920 -2388
rect 1156 -2395 1189 -2387
rect 1614 -2375 1647 -2367
rect 1614 -2392 1622 -2375
rect 1639 -2377 1647 -2375
rect 1883 -2376 1916 -2368
rect 1883 -2377 1891 -2376
rect 1639 -2392 1668 -2377
rect 1710 -2392 1723 -2377
rect 1783 -2392 1796 -2377
rect 1860 -2392 1891 -2377
rect 1614 -2400 1647 -2392
rect 1883 -2393 1891 -2392
rect 1908 -2393 1916 -2376
rect 1883 -2401 1916 -2393
rect 2037 -2376 2070 -2368
rect 2037 -2393 2045 -2376
rect 2062 -2377 2070 -2376
rect 2306 -2375 2339 -2367
rect 2306 -2377 2314 -2375
rect 2062 -2392 2093 -2377
rect 2157 -2392 2170 -2377
rect 2230 -2392 2243 -2377
rect 2285 -2392 2314 -2377
rect 2331 -2392 2339 -2375
rect 2062 -2393 2070 -2392
rect 2037 -2401 2070 -2393
rect 2306 -2400 2339 -2392
rect 2764 -2375 2797 -2367
rect 2764 -2392 2772 -2375
rect 2789 -2377 2797 -2375
rect 3033 -2376 3066 -2368
rect 3033 -2377 3041 -2376
rect 2789 -2392 2818 -2377
rect 2860 -2392 2873 -2377
rect 2933 -2392 2946 -2377
rect 3010 -2392 3041 -2377
rect 2764 -2400 2797 -2392
rect 3033 -2393 3041 -2392
rect 3058 -2393 3066 -2376
rect 3033 -2401 3066 -2393
rect 3187 -2376 3220 -2368
rect 3187 -2393 3195 -2376
rect 3212 -2377 3220 -2376
rect 3456 -2375 3489 -2367
rect 3456 -2377 3464 -2375
rect 3212 -2392 3243 -2377
rect 3307 -2392 3320 -2377
rect 3380 -2392 3393 -2377
rect 3435 -2392 3464 -2377
rect 3481 -2392 3489 -2375
rect 3212 -2393 3220 -2392
rect 3187 -2401 3220 -2393
rect 3456 -2400 3489 -2392
rect 3914 -2375 3947 -2367
rect 3914 -2392 3922 -2375
rect 3939 -2377 3947 -2375
rect 4183 -2376 4216 -2368
rect 4183 -2377 4191 -2376
rect 3939 -2392 3968 -2377
rect 4010 -2392 4023 -2377
rect 4083 -2392 4096 -2377
rect 4160 -2392 4191 -2377
rect 3914 -2400 3947 -2392
rect 4183 -2393 4191 -2392
rect 4208 -2393 4216 -2376
rect 4183 -2401 4216 -2393
rect 4337 -2376 4370 -2368
rect 4337 -2393 4345 -2376
rect 4362 -2377 4370 -2376
rect 4606 -2375 4639 -2367
rect 4606 -2377 4614 -2375
rect 4362 -2392 4393 -2377
rect 4457 -2392 4470 -2377
rect 4530 -2392 4543 -2377
rect 4585 -2392 4614 -2377
rect 4631 -2392 4639 -2375
rect 4362 -2393 4370 -2392
rect 4337 -2401 4370 -2393
rect 4606 -2400 4639 -2392
rect 5064 -2375 5097 -2367
rect 5064 -2392 5072 -2375
rect 5089 -2377 5097 -2375
rect 5333 -2376 5366 -2368
rect 5333 -2377 5341 -2376
rect 5089 -2392 5118 -2377
rect 5160 -2392 5173 -2377
rect 5233 -2392 5246 -2377
rect 5310 -2392 5341 -2377
rect 5064 -2400 5097 -2392
rect 5333 -2393 5341 -2392
rect 5358 -2393 5366 -2376
rect 5333 -2401 5366 -2393
rect 5487 -2376 5520 -2368
rect 5487 -2393 5495 -2376
rect 5512 -2377 5520 -2376
rect 5756 -2375 5789 -2367
rect 5756 -2377 5764 -2375
rect 5512 -2392 5543 -2377
rect 5607 -2392 5620 -2377
rect 5680 -2392 5693 -2377
rect 5735 -2392 5764 -2377
rect 5781 -2392 5789 -2375
rect 5512 -2393 5520 -2392
rect 5487 -2401 5520 -2393
rect 5756 -2400 5789 -2392
rect 6214 -2375 6247 -2367
rect 6214 -2392 6222 -2375
rect 6239 -2377 6247 -2375
rect 6483 -2376 6516 -2368
rect 6483 -2377 6491 -2376
rect 6239 -2392 6268 -2377
rect 6310 -2392 6323 -2377
rect 6383 -2392 6396 -2377
rect 6460 -2392 6491 -2377
rect 6214 -2400 6247 -2392
rect 6483 -2393 6491 -2392
rect 6508 -2393 6516 -2376
rect 6483 -2401 6516 -2393
rect 6637 -2376 6670 -2368
rect 6637 -2393 6645 -2376
rect 6662 -2377 6670 -2376
rect 6906 -2375 6939 -2367
rect 6906 -2377 6914 -2375
rect 6662 -2392 6693 -2377
rect 6757 -2392 6770 -2377
rect 6830 -2392 6843 -2377
rect 6885 -2392 6914 -2377
rect 6931 -2392 6939 -2375
rect 6662 -2393 6670 -2392
rect 6637 -2401 6670 -2393
rect 6906 -2400 6939 -2392
rect 7364 -2375 7397 -2367
rect 7364 -2392 7372 -2375
rect 7389 -2377 7397 -2375
rect 7633 -2376 7666 -2368
rect 7633 -2377 7641 -2376
rect 7389 -2392 7418 -2377
rect 7460 -2392 7473 -2377
rect 7533 -2392 7546 -2377
rect 7610 -2392 7641 -2377
rect 7364 -2400 7397 -2392
rect 7633 -2393 7641 -2392
rect 7658 -2393 7666 -2376
rect 7633 -2401 7666 -2393
rect 7787 -2376 7820 -2368
rect 7787 -2393 7795 -2376
rect 7812 -2377 7820 -2376
rect 8056 -2375 8089 -2367
rect 8056 -2377 8064 -2375
rect 7812 -2392 7843 -2377
rect 7907 -2392 7920 -2377
rect 7980 -2392 7993 -2377
rect 8035 -2392 8064 -2377
rect 8081 -2392 8089 -2375
rect 7812 -2393 7820 -2392
rect 7787 -2401 7820 -2393
rect 8056 -2400 8089 -2392
rect 8514 -2375 8547 -2367
rect 8514 -2392 8522 -2375
rect 8539 -2377 8547 -2375
rect 8783 -2376 8816 -2368
rect 8783 -2377 8791 -2376
rect 8539 -2392 8568 -2377
rect 8610 -2392 8623 -2377
rect 8683 -2392 8696 -2377
rect 8760 -2392 8791 -2377
rect 8514 -2400 8547 -2392
rect 8783 -2393 8791 -2392
rect 8808 -2393 8816 -2376
rect 8783 -2401 8816 -2393
rect 8937 -2376 8970 -2368
rect 8937 -2393 8945 -2376
rect 8962 -2377 8970 -2376
rect 9206 -2375 9239 -2367
rect 9206 -2377 9214 -2375
rect 8962 -2392 8993 -2377
rect 9057 -2392 9070 -2377
rect 9130 -2392 9143 -2377
rect 9185 -2392 9214 -2377
rect 9231 -2392 9239 -2375
rect 8962 -2393 8970 -2392
rect 8937 -2401 8970 -2393
rect 9206 -2400 9239 -2392
<< polycont >>
rect 472 -2389 489 -2372
rect 741 -2388 758 -2371
rect 895 -2388 912 -2371
rect 1164 -2387 1181 -2370
rect 1622 -2392 1639 -2375
rect 1891 -2393 1908 -2376
rect 2045 -2393 2062 -2376
rect 2314 -2392 2331 -2375
rect 2772 -2392 2789 -2375
rect 3041 -2393 3058 -2376
rect 3195 -2393 3212 -2376
rect 3464 -2392 3481 -2375
rect 3922 -2392 3939 -2375
rect 4191 -2393 4208 -2376
rect 4345 -2393 4362 -2376
rect 4614 -2392 4631 -2375
rect 5072 -2392 5089 -2375
rect 5341 -2393 5358 -2376
rect 5495 -2393 5512 -2376
rect 5764 -2392 5781 -2375
rect 6222 -2392 6239 -2375
rect 6491 -2393 6508 -2376
rect 6645 -2393 6662 -2376
rect 6914 -2392 6931 -2375
rect 7372 -2392 7389 -2375
rect 7641 -2393 7658 -2376
rect 7795 -2393 7812 -2376
rect 8064 -2392 8081 -2375
rect 8522 -2392 8539 -2375
rect 8791 -2393 8808 -2376
rect 8945 -2393 8962 -2376
rect 9214 -2392 9231 -2375
<< locali >>
rect 800 -1913 812 -1896
rect 829 -1913 841 -1896
rect 1375 -1913 1387 -1896
rect 1404 -1913 1416 -1896
rect 1950 -1913 1962 -1896
rect 1979 -1913 1991 -1896
rect 2525 -1913 2537 -1896
rect 2554 -1913 2566 -1896
rect 3100 -1913 3112 -1896
rect 3129 -1913 3141 -1896
rect 3675 -1913 3687 -1896
rect 3704 -1913 3716 -1896
rect 4250 -1913 4262 -1896
rect 4279 -1913 4291 -1896
rect 4825 -1913 4837 -1896
rect 4854 -1913 4866 -1896
rect 5400 -1913 5412 -1896
rect 5429 -1913 5441 -1896
rect 5975 -1913 5987 -1896
rect 6004 -1913 6016 -1896
rect 6550 -1913 6562 -1896
rect 6579 -1913 6591 -1896
rect 7125 -1913 7137 -1896
rect 7154 -1913 7166 -1896
rect 7700 -1913 7712 -1896
rect 7729 -1913 7741 -1896
rect 8275 -1913 8287 -1896
rect 8304 -1913 8316 -1896
rect 8850 -1913 8862 -1896
rect 8879 -1913 8891 -1896
rect 9411 -1913 9423 -1896
rect 9440 -1913 9452 -1896
rect 761 -2200 812 -2183
rect 829 -2200 841 -2183
rect 8904 -2184 8940 -2183
rect 1340 -2201 1387 -2184
rect 1404 -2201 1416 -2184
rect 1915 -2201 1962 -2184
rect 1979 -2201 1991 -2184
rect 2490 -2201 2537 -2184
rect 2554 -2201 2566 -2184
rect 3065 -2201 3112 -2184
rect 3129 -2201 3141 -2184
rect 3640 -2201 3687 -2184
rect 3704 -2201 3716 -2184
rect 4215 -2201 4262 -2184
rect 4279 -2201 4291 -2184
rect 4790 -2201 4837 -2184
rect 4854 -2201 4866 -2184
rect 5365 -2201 5412 -2184
rect 5429 -2201 5441 -2184
rect 5940 -2201 5987 -2184
rect 6004 -2201 6016 -2184
rect 6515 -2201 6562 -2184
rect 6579 -2201 6591 -2184
rect 7090 -2201 7137 -2184
rect 7154 -2201 7166 -2184
rect 7665 -2201 7712 -2184
rect 7729 -2201 7741 -2184
rect 8240 -2201 8287 -2184
rect 8304 -2201 8316 -2184
rect 8815 -2201 8862 -2184
rect 8879 -2200 8940 -2184
rect 8879 -2201 8935 -2200
rect 518 -2364 529 -2347
rect 549 -2364 560 -2347
rect 668 -2348 685 -2297
rect 817 -2326 834 -2315
rect 805 -2343 817 -2326
rect 834 -2343 846 -2326
rect 967 -2347 984 -2297
rect 1105 -2345 1122 -2342
rect 464 -2372 497 -2364
rect 646 -2365 668 -2348
rect 685 -2365 710 -2348
rect 464 -2389 472 -2372
rect 489 -2389 497 -2372
rect 733 -2371 766 -2363
rect 733 -2388 741 -2371
rect 758 -2388 766 -2371
rect 464 -2397 497 -2389
rect 531 -2395 548 -2389
rect 472 -2503 489 -2397
rect 518 -2412 531 -2395
rect 548 -2412 669 -2395
rect 686 -2412 710 -2395
rect 733 -2396 766 -2388
rect 887 -2371 920 -2363
rect 943 -2364 967 -2347
rect 984 -2364 1007 -2347
rect 1093 -2364 1104 -2347
rect 1124 -2364 1135 -2347
rect 1681 -2350 1698 -2347
rect 1819 -2352 1836 -2297
rect 1966 -2327 1983 -2316
rect 1954 -2344 1966 -2327
rect 1983 -2344 1995 -2327
rect 2117 -2352 2134 -2297
rect 2255 -2350 2272 -2347
rect 2831 -2350 2848 -2347
rect 2969 -2352 2986 -2297
rect 3109 -2328 3126 -2317
rect 3097 -2345 3109 -2328
rect 3126 -2345 3138 -2328
rect 3267 -2352 3284 -2297
rect 3405 -2350 3422 -2347
rect 3981 -2350 3998 -2347
rect 4119 -2352 4136 -2297
rect 4266 -2329 4283 -2318
rect 4254 -2346 4266 -2329
rect 4283 -2346 4295 -2329
rect 4417 -2352 4434 -2297
rect 4555 -2350 4572 -2347
rect 5131 -2350 5148 -2347
rect 5269 -2352 5286 -2297
rect 5406 -2327 5423 -2316
rect 5394 -2344 5406 -2327
rect 5423 -2344 5435 -2327
rect 5567 -2352 5584 -2297
rect 5705 -2350 5722 -2347
rect 6281 -2350 6298 -2347
rect 6419 -2352 6436 -2297
rect 6574 -2327 6591 -2316
rect 6562 -2344 6574 -2327
rect 6591 -2344 6603 -2327
rect 6717 -2352 6734 -2297
rect 6855 -2350 6872 -2347
rect 7431 -2350 7448 -2347
rect 7569 -2352 7586 -2297
rect 7719 -2327 7736 -2316
rect 7707 -2344 7719 -2327
rect 7736 -2344 7748 -2327
rect 7867 -2352 7884 -2297
rect 8005 -2350 8022 -2347
rect 8581 -2350 8598 -2347
rect 8719 -2352 8736 -2297
rect 8876 -2325 8893 -2314
rect 8864 -2342 8876 -2325
rect 8893 -2342 8905 -2325
rect 9017 -2352 9034 -2297
rect 9155 -2350 9172 -2347
rect 1105 -2370 1122 -2365
rect 1156 -2370 1189 -2362
rect 887 -2388 895 -2371
rect 912 -2388 920 -2371
rect 887 -2396 920 -2388
rect 1156 -2387 1164 -2370
rect 1181 -2387 1189 -2370
rect 531 -2417 548 -2412
rect 669 -2462 686 -2412
rect 741 -2426 758 -2396
rect 741 -2454 758 -2443
rect 896 -2426 913 -2396
rect 943 -2411 968 -2394
rect 985 -2411 1105 -2394
rect 1122 -2411 1135 -2394
rect 1156 -2395 1189 -2387
rect 1614 -2375 1647 -2367
rect 1668 -2369 1679 -2352
rect 1699 -2369 1710 -2352
rect 1796 -2369 1819 -2352
rect 1836 -2369 1860 -2352
rect 1681 -2375 1698 -2370
rect 1614 -2392 1622 -2375
rect 1639 -2392 1647 -2375
rect 896 -2454 913 -2443
rect 968 -2546 985 -2411
rect 1165 -2496 1182 -2395
rect 1614 -2400 1647 -2392
rect 1883 -2376 1916 -2368
rect 1883 -2393 1891 -2376
rect 1908 -2393 1916 -2376
rect 1621 -2495 1638 -2400
rect 1668 -2417 1681 -2400
rect 1698 -2417 1818 -2400
rect 1835 -2417 1860 -2400
rect 1883 -2401 1916 -2393
rect 2037 -2376 2070 -2368
rect 2093 -2369 2117 -2352
rect 2134 -2369 2157 -2352
rect 2243 -2369 2254 -2352
rect 2274 -2369 2285 -2352
rect 2255 -2375 2272 -2370
rect 2306 -2375 2339 -2367
rect 2037 -2393 2045 -2376
rect 2062 -2393 2070 -2376
rect 2037 -2401 2070 -2393
rect 2306 -2392 2314 -2375
rect 2331 -2392 2339 -2375
rect 2306 -2400 2339 -2392
rect 2764 -2375 2797 -2367
rect 2818 -2369 2829 -2352
rect 2849 -2369 2860 -2352
rect 2946 -2369 2969 -2352
rect 2986 -2369 3010 -2352
rect 2831 -2375 2848 -2370
rect 2764 -2392 2772 -2375
rect 2789 -2392 2797 -2375
rect 2764 -2400 2797 -2392
rect 3033 -2376 3066 -2368
rect 3187 -2376 3220 -2368
rect 3243 -2369 3267 -2352
rect 3284 -2369 3307 -2352
rect 3393 -2369 3404 -2352
rect 3424 -2369 3435 -2352
rect 3405 -2375 3422 -2370
rect 3456 -2375 3489 -2367
rect 3033 -2393 3041 -2376
rect 3058 -2393 3083 -2376
rect 3170 -2393 3195 -2376
rect 3212 -2393 3220 -2376
rect 1818 -2609 1835 -2417
rect 1891 -2426 1908 -2401
rect 2046 -2426 2063 -2401
rect 2093 -2417 2118 -2400
rect 2135 -2417 2255 -2400
rect 2272 -2417 2285 -2400
rect 2118 -2684 2135 -2417
rect 2314 -2500 2331 -2400
rect 2773 -2501 2790 -2400
rect 2818 -2417 2831 -2400
rect 2848 -2417 2968 -2400
rect 2985 -2417 3010 -2400
rect 3033 -2401 3066 -2393
rect 3187 -2401 3220 -2393
rect 3456 -2392 3464 -2375
rect 3481 -2392 3489 -2375
rect 3456 -2400 3489 -2392
rect 3914 -2375 3947 -2367
rect 3968 -2369 3979 -2352
rect 3999 -2369 4010 -2352
rect 4096 -2369 4119 -2352
rect 4136 -2369 4160 -2352
rect 3981 -2375 3998 -2370
rect 3914 -2392 3922 -2375
rect 3939 -2392 3947 -2375
rect 3914 -2400 3947 -2392
rect 4183 -2376 4216 -2368
rect 4337 -2376 4370 -2368
rect 4393 -2369 4417 -2352
rect 4434 -2369 4457 -2352
rect 4543 -2369 4554 -2352
rect 4574 -2369 4585 -2352
rect 4555 -2375 4572 -2370
rect 4606 -2375 4639 -2367
rect 4183 -2393 4191 -2376
rect 4208 -2393 4233 -2376
rect 4320 -2393 4345 -2376
rect 4362 -2393 4370 -2376
rect 2968 -2755 2985 -2417
rect 3041 -2426 3058 -2401
rect 3041 -2454 3058 -2443
rect 3195 -2426 3212 -2401
rect 3243 -2418 3268 -2400
rect 3285 -2417 3405 -2400
rect 3422 -2417 3435 -2400
rect 3285 -2418 3307 -2417
rect 3195 -2454 3212 -2443
rect 3268 -2835 3285 -2418
rect 3465 -2499 3482 -2400
rect 3923 -2501 3940 -2400
rect 3968 -2417 3981 -2400
rect 3998 -2417 4118 -2400
rect 4135 -2417 4160 -2400
rect 4183 -2401 4216 -2393
rect 4337 -2401 4370 -2393
rect 4606 -2392 4614 -2375
rect 4631 -2392 4639 -2375
rect 4606 -2400 4639 -2392
rect 5064 -2375 5097 -2367
rect 5118 -2369 5129 -2352
rect 5149 -2369 5160 -2352
rect 5246 -2369 5269 -2352
rect 5286 -2369 5310 -2352
rect 5131 -2375 5148 -2370
rect 5064 -2392 5072 -2375
rect 5089 -2392 5097 -2375
rect 5064 -2400 5097 -2392
rect 5333 -2376 5366 -2368
rect 5487 -2376 5520 -2368
rect 5543 -2369 5567 -2352
rect 5584 -2369 5607 -2352
rect 5693 -2369 5704 -2352
rect 5724 -2369 5735 -2352
rect 5705 -2375 5722 -2370
rect 5756 -2375 5789 -2367
rect 5333 -2393 5341 -2376
rect 5358 -2393 5383 -2376
rect 5470 -2393 5495 -2376
rect 5512 -2393 5520 -2376
rect 4118 -2919 4135 -2417
rect 4188 -2426 4205 -2401
rect 4188 -2454 4205 -2443
rect 4347 -2427 4364 -2401
rect 4393 -2417 4418 -2400
rect 4435 -2417 4555 -2400
rect 4572 -2417 4585 -2400
rect 4347 -2454 4364 -2444
rect 4418 -2990 4435 -2417
rect 4614 -2503 4631 -2400
rect 5072 -2497 5089 -2400
rect 5118 -2417 5131 -2400
rect 5148 -2417 5268 -2400
rect 5285 -2417 5310 -2400
rect 5333 -2401 5366 -2393
rect 5487 -2401 5520 -2393
rect 5756 -2392 5764 -2375
rect 5781 -2392 5789 -2375
rect 5756 -2400 5789 -2392
rect 6214 -2375 6247 -2367
rect 6268 -2369 6279 -2352
rect 6299 -2369 6310 -2352
rect 6396 -2369 6419 -2352
rect 6436 -2369 6460 -2352
rect 6281 -2375 6298 -2370
rect 6214 -2392 6222 -2375
rect 6239 -2392 6247 -2375
rect 6214 -2400 6247 -2392
rect 6483 -2376 6516 -2368
rect 6637 -2376 6670 -2368
rect 6693 -2369 6717 -2352
rect 6734 -2369 6757 -2352
rect 6843 -2369 6854 -2352
rect 6874 -2369 6885 -2352
rect 6855 -2375 6872 -2370
rect 6906 -2375 6939 -2367
rect 6483 -2393 6491 -2376
rect 6508 -2393 6533 -2376
rect 6620 -2393 6645 -2376
rect 6662 -2393 6670 -2376
rect 5268 -3008 5285 -2417
rect 5340 -2426 5357 -2401
rect 5340 -2454 5357 -2443
rect 5495 -2426 5512 -2401
rect 5543 -2417 5568 -2400
rect 5585 -2417 5705 -2400
rect 5722 -2417 5735 -2400
rect 5495 -2454 5512 -2443
rect 5568 -2921 5585 -2417
rect 5765 -2499 5782 -2400
rect 6222 -2495 6239 -2400
rect 6268 -2417 6281 -2400
rect 6298 -2417 6418 -2400
rect 6435 -2417 6460 -2400
rect 6483 -2401 6516 -2393
rect 6637 -2401 6670 -2393
rect 6906 -2392 6914 -2375
rect 6931 -2392 6939 -2375
rect 6906 -2400 6939 -2392
rect 7364 -2375 7397 -2367
rect 7418 -2369 7429 -2352
rect 7449 -2369 7460 -2352
rect 7546 -2369 7569 -2352
rect 7586 -2369 7610 -2352
rect 7431 -2375 7448 -2370
rect 7364 -2392 7372 -2375
rect 7389 -2392 7397 -2375
rect 7364 -2400 7397 -2392
rect 7633 -2376 7666 -2368
rect 7787 -2376 7820 -2368
rect 7843 -2369 7867 -2352
rect 7884 -2369 7907 -2352
rect 7993 -2369 8004 -2352
rect 8024 -2369 8035 -2352
rect 8005 -2375 8022 -2370
rect 8056 -2375 8089 -2367
rect 7633 -2393 7641 -2376
rect 7658 -2393 7683 -2376
rect 7770 -2393 7795 -2376
rect 7812 -2393 7820 -2376
rect 6418 -2841 6435 -2417
rect 6491 -2427 6508 -2401
rect 6491 -2454 6508 -2444
rect 6644 -2427 6661 -2401
rect 6693 -2417 6718 -2400
rect 6735 -2417 6855 -2400
rect 6872 -2417 6885 -2400
rect 6644 -2454 6661 -2444
rect 6718 -2769 6735 -2417
rect 6914 -2499 6931 -2400
rect 7372 -2499 7389 -2400
rect 7418 -2417 7431 -2400
rect 7448 -2417 7568 -2400
rect 7585 -2417 7610 -2400
rect 7633 -2401 7666 -2393
rect 7787 -2401 7820 -2393
rect 8056 -2392 8064 -2375
rect 8081 -2392 8089 -2375
rect 8056 -2400 8089 -2392
rect 8514 -2375 8547 -2367
rect 8568 -2369 8579 -2352
rect 8599 -2369 8610 -2352
rect 8696 -2369 8719 -2352
rect 8736 -2369 8760 -2352
rect 8581 -2375 8598 -2370
rect 8514 -2392 8522 -2375
rect 8539 -2392 8547 -2375
rect 8514 -2400 8547 -2392
rect 8783 -2376 8816 -2368
rect 8937 -2376 8970 -2368
rect 8993 -2369 9017 -2352
rect 9034 -2369 9057 -2352
rect 9143 -2369 9154 -2352
rect 9174 -2369 9185 -2352
rect 9155 -2375 9172 -2370
rect 9206 -2375 9239 -2367
rect 8783 -2393 8791 -2376
rect 8808 -2393 8833 -2376
rect 8920 -2393 8945 -2376
rect 8962 -2393 8970 -2376
rect 7568 -2706 7585 -2417
rect 7642 -2426 7659 -2401
rect 7642 -2454 7659 -2443
rect 7795 -2426 7812 -2401
rect 7843 -2417 7868 -2400
rect 7885 -2417 8005 -2400
rect 8022 -2417 8035 -2400
rect 7795 -2454 7812 -2443
rect 7868 -2643 7885 -2417
rect 8064 -2502 8081 -2400
rect 8522 -2500 8539 -2400
rect 8568 -2417 8581 -2400
rect 8598 -2417 8718 -2400
rect 8735 -2417 8760 -2400
rect 8783 -2401 8816 -2393
rect 8937 -2401 8970 -2393
rect 9206 -2392 9214 -2375
rect 9231 -2392 9239 -2375
rect 9206 -2400 9239 -2392
rect 8718 -2593 8735 -2417
rect 8791 -2425 8808 -2401
rect 8791 -2454 8808 -2442
rect 8943 -2426 8960 -2401
rect 8993 -2417 9018 -2400
rect 9035 -2417 9155 -2400
rect 9172 -2417 9185 -2400
rect 8943 -2454 8960 -2443
rect 9018 -2543 9035 -2417
rect 9216 -2487 9233 -2400
rect 9206 -2494 9236 -2487
rect 9206 -2518 9209 -2494
rect 9233 -2518 9236 -2494
rect 9206 -2521 9236 -2518
rect -3215 -4451 -3198 -4417
rect -2065 -4450 -2048 -4417
rect -883 -4450 -866 -4417
rect 298 -4450 315 -4417
rect 1479 -4450 1496 -4417
rect 2661 -4450 2678 -4417
rect 3843 -4450 3860 -4417
rect 5025 -4450 5042 -4417
rect 6207 -4450 6224 -4417
rect 7389 -4450 7406 -4417
rect 8571 -4450 8588 -4417
rect 9755 -4450 9772 -4417
rect 10939 -4450 10956 -4417
rect 12126 -4450 12143 -4417
rect 13313 -4450 13330 -4417
rect 14196 -4434 14231 -4417
rect 14214 -4450 14231 -4434
rect -3215 -4589 -3198 -4557
rect -2065 -4589 -2048 -4556
rect -883 -4542 -866 -4539
rect -883 -4589 -866 -4559
rect 298 -4589 315 -4556
rect 1479 -4589 1496 -4556
rect 2661 -4589 2678 -4556
rect 3843 -4589 3860 -4556
rect 5025 -4589 5042 -4556
rect 6207 -4589 6224 -4556
rect 7389 -4589 7406 -4556
rect 8571 -4589 8588 -4556
rect 9755 -4589 9772 -4556
rect 10939 -4589 10956 -4557
rect 12126 -4589 12143 -4556
rect 13313 -4589 13330 -4556
rect 14214 -4572 14231 -4556
rect 14179 -4589 14231 -4572
rect -3215 -7177 -3198 -7152
rect -2065 -7176 -2048 -7152
rect -883 -7176 -866 -7152
rect 298 -7176 315 -7152
rect 1479 -7176 1496 -7152
rect 2661 -7176 2678 -7152
rect 3843 -7176 3860 -7152
rect 5025 -7176 5042 -7152
rect 6207 -7176 6224 -7152
rect 7389 -7176 7406 -7152
rect 8571 -7176 8588 -7152
rect 9755 -7176 9772 -7152
rect 10939 -7176 10956 -7152
rect 12126 -7176 12143 -7152
rect 13313 -7176 13330 -7152
rect 14196 -7169 14231 -7152
rect 14214 -7176 14231 -7169
rect -3215 -7321 -3198 -7291
rect -2065 -7321 -2048 -7290
rect -883 -7321 -866 -7290
rect 298 -7321 315 -7290
rect 1479 -7321 1496 -7290
rect 2661 -7321 2678 -7290
rect 3843 -7321 3860 -7290
rect 5025 -7321 5042 -7290
rect 6207 -7321 6224 -7290
rect 7389 -7321 7406 -7290
rect 8571 -7321 8588 -7290
rect 9755 -7321 9772 -7290
rect 10939 -7321 10956 -7290
rect 12126 -7321 12143 -7290
rect 13313 -7321 13330 -7290
rect 14214 -7304 14231 -7290
rect 14196 -7321 14231 -7304
<< viali >>
rect 601 -1408 618 -1391
rect 1176 -1409 1193 -1392
rect 1751 -1411 1768 -1394
rect 2326 -1411 2343 -1394
rect 2901 -1409 2918 -1392
rect 3476 -1406 3493 -1389
rect 4051 -1404 4068 -1387
rect 4626 -1404 4643 -1387
rect 5201 -1409 5218 -1392
rect 5776 -1406 5793 -1389
rect 6351 -1410 6368 -1393
rect 6926 -1411 6943 -1394
rect 7501 -1407 7518 -1390
rect 8076 -1411 8093 -1394
rect 8651 -1407 8668 -1390
rect 9226 -1408 9243 -1391
rect 812 -1913 829 -1896
rect 1387 -1913 1404 -1896
rect 1962 -1913 1979 -1896
rect 2537 -1913 2554 -1896
rect 3112 -1913 3129 -1896
rect 3687 -1913 3704 -1896
rect 4262 -1913 4279 -1896
rect 4837 -1913 4854 -1896
rect 5412 -1913 5429 -1896
rect 5987 -1913 6004 -1896
rect 6562 -1913 6579 -1896
rect 7137 -1913 7154 -1896
rect 7712 -1913 7729 -1896
rect 8287 -1913 8304 -1896
rect 8862 -1913 8879 -1896
rect 9423 -1913 9440 -1896
rect 668 -2297 685 -2280
rect 529 -2347 549 -2344
rect 529 -2364 531 -2347
rect 531 -2364 548 -2347
rect 548 -2364 549 -2347
rect 967 -2297 984 -2280
rect 817 -2343 834 -2327
rect 817 -2344 834 -2343
rect 1819 -2297 1836 -2280
rect 1104 -2347 1124 -2345
rect 1104 -2364 1105 -2347
rect 1105 -2364 1122 -2347
rect 1122 -2364 1124 -2347
rect 1679 -2352 1699 -2350
rect 2117 -2297 2134 -2280
rect 1966 -2344 1983 -2328
rect 1966 -2345 1983 -2344
rect 2969 -2297 2986 -2280
rect 2254 -2352 2274 -2350
rect 2829 -2352 2849 -2350
rect 3267 -2297 3284 -2280
rect 3109 -2345 3126 -2329
rect 3109 -2346 3126 -2345
rect 4119 -2297 4136 -2280
rect 3404 -2352 3424 -2350
rect 3979 -2352 3999 -2350
rect 4417 -2297 4434 -2280
rect 4266 -2346 4283 -2330
rect 4266 -2347 4283 -2346
rect 5269 -2297 5286 -2280
rect 4554 -2352 4574 -2350
rect 5129 -2352 5149 -2350
rect 5567 -2297 5584 -2280
rect 5406 -2344 5423 -2328
rect 5406 -2345 5423 -2344
rect 6419 -2297 6436 -2280
rect 5704 -2352 5724 -2350
rect 6279 -2352 6299 -2350
rect 6717 -2297 6734 -2280
rect 6574 -2344 6591 -2328
rect 6574 -2345 6591 -2344
rect 7569 -2297 7586 -2280
rect 6854 -2352 6874 -2350
rect 7429 -2352 7449 -2350
rect 7867 -2297 7884 -2280
rect 7719 -2344 7736 -2328
rect 7719 -2345 7736 -2344
rect 8719 -2297 8736 -2280
rect 8004 -2352 8024 -2350
rect 8579 -2352 8599 -2350
rect 9017 -2297 9034 -2280
rect 8876 -2342 8893 -2326
rect 8876 -2343 8893 -2342
rect 9154 -2352 9174 -2350
rect 1104 -2365 1124 -2364
rect 741 -2443 758 -2426
rect 1679 -2369 1681 -2352
rect 1681 -2369 1698 -2352
rect 1698 -2369 1699 -2352
rect 1679 -2370 1699 -2369
rect 896 -2443 913 -2426
rect 669 -2479 686 -2462
rect 472 -2520 489 -2503
rect 1165 -2513 1182 -2496
rect 2254 -2369 2255 -2352
rect 2255 -2369 2272 -2352
rect 2272 -2369 2274 -2352
rect 2254 -2370 2274 -2369
rect 2829 -2369 2831 -2352
rect 2831 -2369 2848 -2352
rect 2848 -2369 2849 -2352
rect 2829 -2370 2849 -2369
rect 3404 -2369 3405 -2352
rect 3405 -2369 3422 -2352
rect 3422 -2369 3424 -2352
rect 3404 -2370 3424 -2369
rect 1621 -2512 1638 -2495
rect 968 -2563 985 -2546
rect 1891 -2443 1908 -2426
rect 2046 -2443 2063 -2426
rect 1818 -2626 1835 -2609
rect 2314 -2517 2331 -2500
rect 3979 -2369 3981 -2352
rect 3981 -2369 3998 -2352
rect 3998 -2369 3999 -2352
rect 3979 -2370 3999 -2369
rect 4554 -2369 4555 -2352
rect 4555 -2369 4572 -2352
rect 4572 -2369 4574 -2352
rect 4554 -2370 4574 -2369
rect 2773 -2518 2790 -2501
rect 2118 -2701 2135 -2684
rect 3041 -2443 3058 -2426
rect 3195 -2443 3212 -2426
rect 2968 -2772 2985 -2755
rect 3465 -2516 3482 -2499
rect 5129 -2369 5131 -2352
rect 5131 -2369 5148 -2352
rect 5148 -2369 5149 -2352
rect 5129 -2370 5149 -2369
rect 5704 -2369 5705 -2352
rect 5705 -2369 5722 -2352
rect 5722 -2369 5724 -2352
rect 5704 -2370 5724 -2369
rect 3923 -2518 3940 -2501
rect 3268 -2852 3285 -2835
rect 4188 -2443 4205 -2426
rect 4347 -2444 4364 -2427
rect 4118 -2936 4135 -2919
rect 4614 -2520 4631 -2503
rect 6279 -2369 6281 -2352
rect 6281 -2369 6298 -2352
rect 6298 -2369 6299 -2352
rect 6279 -2370 6299 -2369
rect 6854 -2369 6855 -2352
rect 6855 -2369 6872 -2352
rect 6872 -2369 6874 -2352
rect 6854 -2370 6874 -2369
rect 5072 -2514 5089 -2497
rect 4418 -3007 4435 -2990
rect 5340 -2443 5357 -2426
rect 5495 -2443 5512 -2426
rect 5765 -2516 5782 -2499
rect 7429 -2369 7431 -2352
rect 7431 -2369 7448 -2352
rect 7448 -2369 7449 -2352
rect 7429 -2370 7449 -2369
rect 8004 -2369 8005 -2352
rect 8005 -2369 8022 -2352
rect 8022 -2369 8024 -2352
rect 8004 -2370 8024 -2369
rect 6222 -2512 6239 -2495
rect 6491 -2444 6508 -2427
rect 6644 -2444 6661 -2427
rect 6914 -2516 6931 -2499
rect 8579 -2369 8581 -2352
rect 8581 -2369 8598 -2352
rect 8598 -2369 8599 -2352
rect 8579 -2370 8599 -2369
rect 9154 -2369 9155 -2352
rect 9155 -2369 9172 -2352
rect 9172 -2369 9174 -2352
rect 9154 -2370 9174 -2369
rect 7372 -2516 7389 -2499
rect 7642 -2443 7659 -2426
rect 7795 -2443 7812 -2426
rect 8064 -2519 8081 -2502
rect 8522 -2517 8539 -2500
rect 8791 -2442 8808 -2425
rect 8943 -2443 8960 -2426
rect 9209 -2518 9233 -2494
rect 9018 -2560 9035 -2543
rect 8718 -2610 8735 -2593
rect 7868 -2660 7885 -2643
rect 7568 -2723 7585 -2706
rect 6718 -2786 6735 -2769
rect 6418 -2858 6435 -2841
rect 5568 -2938 5585 -2921
rect 5268 -3025 5285 -3008
rect -3654 -3606 -3637 -3589
rect -2481 -3606 -2464 -3589
rect -1309 -3606 -1292 -3589
rect -128 -3606 -111 -3589
rect 1058 -3606 1075 -3589
rect 2242 -3606 2259 -3589
rect 3410 -3606 3427 -3589
rect 4599 -3606 4616 -3589
rect 5777 -3606 5794 -3589
rect 6966 -3606 6983 -3589
rect 8132 -3606 8149 -3589
rect 9334 -3606 9351 -3589
rect 10507 -3606 10524 -3589
rect 11679 -3606 11696 -3589
rect 12895 -3606 12912 -3589
rect 13797 -3606 13814 -3589
rect -3215 -4468 -3198 -4451
rect -2065 -4467 -2048 -4450
rect -883 -4467 -866 -4450
rect 298 -4467 315 -4450
rect 1479 -4467 1496 -4450
rect 2661 -4467 2678 -4450
rect 3843 -4467 3860 -4450
rect 5025 -4467 5042 -4450
rect 6207 -4467 6224 -4450
rect 7389 -4467 7406 -4450
rect 8571 -4467 8588 -4450
rect 9755 -4467 9772 -4450
rect 10939 -4467 10956 -4450
rect 12126 -4467 12143 -4450
rect 13313 -4467 13330 -4450
rect 14214 -4467 14231 -4450
rect -3215 -4557 -3198 -4540
rect -2065 -4556 -2048 -4539
rect -883 -4559 -866 -4542
rect 298 -4556 315 -4539
rect 1479 -4556 1496 -4539
rect 2661 -4556 2678 -4539
rect 3843 -4556 3860 -4539
rect 5025 -4556 5042 -4539
rect 6207 -4556 6224 -4539
rect 7389 -4556 7406 -4539
rect 8571 -4556 8588 -4539
rect 9755 -4556 9772 -4539
rect 10939 -4557 10956 -4540
rect 12126 -4556 12143 -4539
rect 13313 -4556 13330 -4539
rect 14214 -4556 14231 -4539
rect -3632 -5418 -3615 -5401
rect -2501 -5419 -2484 -5402
rect -1320 -5419 -1303 -5402
rect -148 -5419 -131 -5402
rect 1030 -5419 1047 -5402
rect 2218 -5419 2235 -5402
rect 3409 -5419 3426 -5402
rect 4591 -5419 4608 -5402
rect 5760 -5419 5777 -5402
rect 6948 -5419 6965 -5402
rect 8127 -5419 8144 -5402
rect 9315 -5419 9332 -5402
rect 10492 -5419 10509 -5402
rect 11670 -5419 11687 -5402
rect 12851 -5419 12868 -5402
rect 13778 -5419 13795 -5402
rect -3634 -6339 -3617 -6322
rect -2486 -6339 -2469 -6322
rect -1305 -6339 -1288 -6322
rect -130 -6339 -113 -6322
rect 1058 -6339 1075 -6322
rect 2242 -6339 2259 -6322
rect 3413 -6339 3430 -6322
rect 4600 -6339 4617 -6322
rect 5788 -6339 5805 -6322
rect 6955 -6339 6972 -6322
rect 8137 -6339 8154 -6322
rect 9323 -6339 9340 -6322
rect 10499 -6339 10516 -6322
rect 11678 -6339 11695 -6322
rect 12880 -6339 12897 -6322
rect 13779 -6339 13796 -6322
rect -3215 -7194 -3198 -7177
rect -2065 -7193 -2048 -7176
rect -883 -7193 -866 -7176
rect 298 -7193 315 -7176
rect 1479 -7193 1496 -7176
rect 2661 -7193 2678 -7176
rect 3843 -7193 3860 -7176
rect 5025 -7193 5042 -7176
rect 6207 -7193 6224 -7176
rect 7389 -7193 7406 -7176
rect 8571 -7193 8588 -7176
rect 9755 -7193 9772 -7176
rect 10939 -7193 10956 -7176
rect 12126 -7193 12143 -7176
rect 13313 -7193 13330 -7176
rect 14214 -7193 14231 -7176
rect -3215 -7291 -3198 -7274
rect -2065 -7290 -2048 -7273
rect -883 -7290 -866 -7273
rect 298 -7290 315 -7273
rect 1479 -7290 1496 -7273
rect 2661 -7290 2678 -7273
rect 3843 -7290 3860 -7273
rect 5025 -7290 5042 -7273
rect 6207 -7290 6224 -7273
rect 7389 -7290 7406 -7273
rect 8571 -7290 8588 -7273
rect 9755 -7290 9772 -7273
rect 10939 -7290 10956 -7273
rect 12126 -7290 12143 -7273
rect 13313 -7290 13330 -7273
rect 14214 -7290 14231 -7273
rect -3643 -8152 -3626 -8135
rect -2508 -8152 -2491 -8135
rect -1333 -8152 -1316 -8135
rect -151 -8152 -134 -8135
rect 1031 -8152 1048 -8135
rect 2213 -8152 2230 -8135
rect 3407 -8152 3424 -8135
rect 4584 -8152 4601 -8135
rect 5767 -8152 5784 -8135
rect 6940 -8152 6957 -8135
rect 8123 -8152 8140 -8135
rect 9306 -8152 9323 -8135
rect 10484 -8152 10501 -8135
rect 11678 -8152 11695 -8135
rect 12873 -8152 12890 -8135
rect 13778 -8152 13795 -8135
<< metal1 >>
rect 519 5034 559 5074
rect 1095 5034 1135 5074
rect 1670 5034 1710 5074
rect 2243 5034 2283 5074
rect 2819 5034 2859 5074
rect 3393 5034 3433 5074
rect 3968 5034 4008 5074
rect 4543 5034 4583 5074
rect 5118 5034 5158 5074
rect 5694 5034 5734 5074
rect 6269 5033 6309 5073
rect 6843 5034 6883 5074
rect 7418 5034 7458 5074
rect 7993 5034 8033 5074
rect 8567 5034 8607 5074
rect 9142 5034 9182 5074
rect -4549 5000 239 5014
rect 126 4838 129 4864
rect 155 4858 158 4864
rect 155 4844 242 4858
rect 155 4838 158 4844
rect 125 4781 157 4784
rect 125 4755 128 4781
rect 154 4775 157 4781
rect 154 4761 239 4775
rect 154 4755 157 4761
rect 125 4752 157 4755
rect -4549 4721 251 4735
rect 127 4695 159 4698
rect 127 4669 130 4695
rect 156 4694 159 4695
rect 156 4680 242 4694
rect 156 4669 159 4680
rect 127 4666 159 4669
rect 125 4597 128 4623
rect 154 4617 157 4623
rect 154 4603 239 4617
rect 154 4597 157 4603
rect 126 4538 158 4541
rect 126 4512 129 4538
rect 155 4534 158 4538
rect 155 4520 240 4534
rect 155 4512 158 4520
rect 126 4509 158 4512
rect -4549 4480 239 4494
rect 126 4458 158 4461
rect 126 4432 129 4458
rect 155 4453 158 4458
rect 155 4439 249 4453
rect 155 4432 158 4439
rect 126 4429 158 4432
rect 125 4356 128 4382
rect 154 4376 157 4382
rect 154 4362 239 4376
rect 154 4356 157 4362
rect 127 4245 159 4248
rect 127 4219 130 4245
rect 156 4237 159 4245
rect 156 4223 239 4237
rect 156 4219 159 4223
rect 127 4216 159 4219
rect -4549 4183 240 4197
rect 127 4159 159 4162
rect 127 4133 130 4159
rect 156 4156 159 4159
rect 156 4142 244 4156
rect 156 4133 159 4142
rect 127 4130 159 4133
rect 125 4059 128 4085
rect 154 4079 157 4085
rect 154 4065 239 4079
rect 154 4059 157 4065
rect 127 4002 159 4005
rect 127 3976 130 4002
rect 156 3996 159 4002
rect 156 3982 239 3996
rect 156 3976 159 3982
rect 127 3973 159 3976
rect -4549 3942 244 3956
rect 127 3918 159 3921
rect 127 3892 130 3918
rect 156 3915 159 3918
rect 156 3901 242 3915
rect 156 3892 159 3901
rect 127 3889 159 3892
rect 126 3818 129 3844
rect 155 3838 158 3844
rect 155 3824 225 3838
rect 231 3824 239 3838
rect 155 3818 158 3824
rect -4549 3741 239 3755
rect -4549 3701 239 3715
rect -4549 3660 239 3674
rect 126 3577 129 3603
rect 155 3597 158 3603
rect 155 3583 247 3597
rect 155 3577 158 3583
rect -4549 3500 240 3514
rect -4549 3460 244 3474
rect -4549 3419 239 3433
rect 126 3336 129 3362
rect 155 3356 158 3362
rect 155 3342 239 3356
rect 155 3336 158 3342
rect -4549 3259 239 3273
rect -4549 3219 243 3233
rect -4549 3178 241 3192
rect 126 3095 129 3121
rect 155 3115 158 3121
rect 155 3101 239 3115
rect 155 3095 158 3101
rect -4549 3018 239 3032
rect -4549 2978 242 2992
rect -4549 2937 239 2951
rect 126 2854 129 2880
rect 155 2874 158 2880
rect 155 2860 239 2874
rect 155 2854 158 2860
rect -4549 2737 239 2751
rect -4549 2697 240 2711
rect -4549 2656 239 2670
rect 125 2573 128 2599
rect 154 2593 157 2599
rect 154 2579 239 2593
rect 154 2573 157 2579
rect -4549 2496 239 2510
rect -4549 2456 239 2470
rect -4549 2415 239 2429
rect 126 2332 129 2358
rect 155 2352 158 2358
rect 155 2338 240 2352
rect 155 2332 158 2338
rect -4549 2255 239 2269
rect -4549 2215 239 2229
rect -4549 2174 239 2188
rect 126 2091 129 2117
rect 155 2111 158 2117
rect 155 2097 239 2111
rect 155 2091 158 2097
rect -4549 2014 239 2028
rect -4549 1974 239 1988
rect -4549 1933 239 1947
rect 126 1850 129 1876
rect 155 1870 158 1876
rect 155 1856 239 1870
rect 155 1850 158 1856
rect -4549 1773 239 1787
rect -4549 1733 241 1747
rect -4549 1692 239 1706
rect 126 1609 129 1635
rect 155 1629 158 1635
rect 155 1615 239 1629
rect 155 1609 158 1615
rect -4549 1532 239 1546
rect -4549 1492 240 1506
rect -4549 1451 244 1465
rect 126 1368 129 1394
rect 155 1388 158 1394
rect 155 1374 251 1388
rect 155 1368 158 1374
rect -4549 1291 239 1305
rect -4549 1251 240 1265
rect -4549 1210 239 1224
rect 125 1127 128 1153
rect 154 1147 157 1153
rect 154 1133 240 1147
rect 154 1127 157 1133
rect -4549 1050 239 1064
rect -4549 1010 242 1024
rect -4549 969 240 983
rect 126 886 129 912
rect 155 906 158 912
rect 155 892 247 906
rect 155 886 158 892
rect -4549 768 239 782
rect -4549 728 242 742
rect -4549 687 239 701
rect 125 604 128 630
rect 154 624 157 630
rect 154 610 239 624
rect 154 604 157 610
rect -4549 527 239 541
rect -4549 487 239 501
rect -4549 446 239 460
rect 127 363 130 389
rect 156 383 159 389
rect 156 369 242 383
rect 156 363 159 369
rect -4549 286 239 300
rect -4549 246 240 260
rect -4549 205 242 219
rect 126 122 129 148
rect 155 142 158 148
rect 155 128 239 142
rect 155 122 158 128
rect -4549 45 239 59
rect -4549 5 239 19
rect -4549 -36 239 -22
rect 126 -93 158 -90
rect 126 -119 129 -93
rect 155 -99 158 -93
rect 155 -113 250 -99
rect 155 -119 158 -113
rect 126 -122 158 -119
rect 126 -178 158 -175
rect 126 -204 129 -178
rect 155 -182 158 -178
rect 155 -196 239 -182
rect 155 -204 158 -196
rect 126 -207 158 -204
rect -4549 -236 246 -222
rect 126 -257 158 -254
rect 126 -283 129 -257
rect 155 -263 158 -257
rect 155 -277 239 -263
rect 155 -283 158 -277
rect 126 -286 158 -283
rect 129 -334 155 -331
rect 155 -354 242 -340
rect 129 -363 155 -360
rect 126 -416 158 -413
rect 126 -442 129 -416
rect 155 -423 158 -416
rect 155 -437 239 -423
rect 155 -442 158 -437
rect 126 -445 158 -442
rect -4549 -477 239 -463
rect 127 -495 159 -492
rect 127 -521 130 -495
rect 156 -504 159 -495
rect 156 -518 239 -504
rect 156 -521 159 -518
rect 127 -524 159 -521
rect 126 -601 129 -575
rect 155 -581 158 -575
rect 155 -595 239 -581
rect 155 -601 158 -595
rect 126 -718 158 -715
rect 126 -744 129 -718
rect 155 -723 158 -718
rect 155 -737 239 -723
rect 155 -744 158 -737
rect 126 -747 158 -744
rect -4549 -777 239 -763
rect 126 -798 158 -795
rect 126 -824 129 -798
rect 155 -804 158 -798
rect 155 -818 239 -804
rect 155 -824 158 -818
rect 126 -827 158 -824
rect 126 -875 158 -872
rect 126 -901 129 -875
rect 155 -881 158 -875
rect 155 -895 239 -881
rect 155 -901 158 -895
rect 126 -904 158 -901
rect 126 -955 158 -952
rect 126 -981 129 -955
rect 155 -964 158 -955
rect 155 -978 241 -964
rect 155 -981 158 -978
rect 126 -984 158 -981
rect -4549 -1018 239 -1004
rect 127 -1042 159 -1039
rect 127 -1068 130 -1042
rect 156 -1045 159 -1042
rect 156 -1059 241 -1045
rect 156 -1068 159 -1059
rect 127 -1071 159 -1068
rect 126 -1142 129 -1116
rect 155 -1122 158 -1116
rect 155 -1136 239 -1122
rect 155 -1142 158 -1136
rect 594 -1386 626 -1383
rect 3469 -1384 3501 -1381
rect 594 -1412 597 -1386
rect 623 -1412 626 -1386
rect 594 -1415 626 -1412
rect 1169 -1387 1201 -1384
rect 1169 -1413 1172 -1387
rect 1198 -1413 1201 -1387
rect 1169 -1416 1201 -1413
rect 1744 -1389 1776 -1386
rect 1744 -1415 1747 -1389
rect 1773 -1415 1776 -1389
rect 1744 -1418 1776 -1415
rect 2319 -1389 2351 -1386
rect 2319 -1415 2322 -1389
rect 2348 -1415 2351 -1389
rect 2319 -1418 2351 -1415
rect 2894 -1387 2926 -1384
rect 2894 -1413 2897 -1387
rect 2923 -1413 2926 -1387
rect 3469 -1410 3472 -1384
rect 3498 -1410 3501 -1384
rect 3469 -1413 3501 -1410
rect 4040 -1382 4080 -1375
rect 4040 -1408 4047 -1382
rect 4073 -1408 4080 -1382
rect 2894 -1416 2926 -1413
rect 4040 -1415 4080 -1408
rect 4619 -1382 4651 -1379
rect 4619 -1408 4622 -1382
rect 4648 -1408 4651 -1382
rect 5769 -1384 5801 -1381
rect 4619 -1411 4651 -1408
rect 5194 -1387 5226 -1384
rect 5194 -1413 5197 -1387
rect 5223 -1413 5226 -1387
rect 5769 -1410 5772 -1384
rect 5798 -1410 5801 -1384
rect 7494 -1385 7526 -1382
rect 5769 -1413 5801 -1410
rect 6344 -1388 6376 -1385
rect 5194 -1416 5226 -1413
rect 6344 -1414 6347 -1388
rect 6373 -1414 6376 -1388
rect 6344 -1417 6376 -1414
rect 6919 -1389 6951 -1386
rect 6919 -1415 6922 -1389
rect 6948 -1415 6951 -1389
rect 7494 -1411 7497 -1385
rect 7523 -1411 7526 -1385
rect 8644 -1385 8676 -1382
rect 7494 -1414 7526 -1411
rect 8069 -1389 8101 -1386
rect 6919 -1418 6951 -1415
rect 8069 -1415 8072 -1389
rect 8098 -1415 8101 -1389
rect 8644 -1411 8647 -1385
rect 8673 -1411 8676 -1385
rect 8644 -1414 8676 -1411
rect 9219 -1386 9251 -1383
rect 9219 -1412 9222 -1386
rect 9248 -1412 9251 -1386
rect 9219 -1415 9251 -1412
rect 8069 -1418 8101 -1415
rect -4549 -1866 242 -1852
rect 126 -1919 129 -1893
rect 155 -1899 158 -1893
rect 806 -1896 835 -1890
rect 155 -1913 239 -1899
rect 806 -1913 812 -1896
rect 829 -1913 835 -1896
rect 1381 -1896 1410 -1890
rect 1381 -1898 1387 -1896
rect 1375 -1912 1387 -1898
rect 155 -1919 158 -1913
rect 806 -1919 835 -1913
rect 1381 -1913 1387 -1912
rect 1404 -1898 1410 -1896
rect 1956 -1896 1985 -1890
rect 1956 -1898 1962 -1896
rect 1404 -1912 1416 -1898
rect 1950 -1912 1962 -1898
rect 1404 -1913 1410 -1912
rect 1381 -1919 1410 -1913
rect 1956 -1913 1962 -1912
rect 1979 -1898 1985 -1896
rect 2531 -1896 2560 -1890
rect 2531 -1898 2537 -1896
rect 1979 -1912 1991 -1898
rect 2525 -1912 2537 -1898
rect 1979 -1913 1985 -1912
rect 1956 -1919 1985 -1913
rect 2531 -1913 2537 -1912
rect 2554 -1898 2560 -1896
rect 3106 -1896 3135 -1890
rect 3106 -1898 3112 -1896
rect 2554 -1912 2566 -1898
rect 3100 -1912 3112 -1898
rect 2554 -1913 2560 -1912
rect 2531 -1919 2560 -1913
rect 3106 -1913 3112 -1912
rect 3129 -1898 3135 -1896
rect 3681 -1896 3710 -1890
rect 3681 -1898 3687 -1896
rect 3129 -1912 3141 -1898
rect 3675 -1912 3687 -1898
rect 3129 -1913 3135 -1912
rect 3106 -1919 3135 -1913
rect 3681 -1913 3687 -1912
rect 3704 -1898 3710 -1896
rect 4256 -1896 4285 -1890
rect 4256 -1898 4262 -1896
rect 3704 -1912 3716 -1898
rect 4250 -1912 4262 -1898
rect 3704 -1913 3710 -1912
rect 3681 -1919 3710 -1913
rect 4256 -1913 4262 -1912
rect 4279 -1898 4285 -1896
rect 4831 -1896 4860 -1890
rect 4831 -1898 4837 -1896
rect 4279 -1912 4291 -1898
rect 4825 -1912 4837 -1898
rect 4279 -1913 4285 -1912
rect 4256 -1919 4285 -1913
rect 4831 -1913 4837 -1912
rect 4854 -1898 4860 -1896
rect 5406 -1896 5435 -1890
rect 5406 -1898 5412 -1896
rect 4854 -1912 4866 -1898
rect 5400 -1912 5412 -1898
rect 4854 -1913 4860 -1912
rect 4831 -1919 4860 -1913
rect 5406 -1913 5412 -1912
rect 5429 -1898 5435 -1896
rect 5981 -1896 6010 -1890
rect 5981 -1898 5987 -1896
rect 5429 -1912 5441 -1898
rect 5975 -1912 5987 -1898
rect 5429 -1913 5435 -1912
rect 5406 -1919 5435 -1913
rect 5981 -1913 5987 -1912
rect 6004 -1898 6010 -1896
rect 6556 -1896 6585 -1890
rect 6556 -1898 6562 -1896
rect 6004 -1912 6016 -1898
rect 6550 -1912 6562 -1898
rect 6004 -1913 6010 -1912
rect 5981 -1919 6010 -1913
rect 6556 -1913 6562 -1912
rect 6579 -1898 6585 -1896
rect 7131 -1896 7160 -1890
rect 7131 -1898 7137 -1896
rect 6579 -1912 6591 -1898
rect 7125 -1912 7137 -1898
rect 6579 -1913 6585 -1912
rect 6556 -1919 6585 -1913
rect 7131 -1913 7137 -1912
rect 7154 -1898 7160 -1896
rect 7706 -1896 7735 -1890
rect 7706 -1898 7712 -1896
rect 7154 -1912 7166 -1898
rect 7700 -1912 7712 -1898
rect 7154 -1913 7160 -1912
rect 7131 -1919 7160 -1913
rect 7706 -1913 7712 -1912
rect 7729 -1898 7735 -1896
rect 8281 -1896 8310 -1890
rect 8281 -1898 8287 -1896
rect 7729 -1912 7741 -1898
rect 8275 -1912 8287 -1898
rect 7729 -1913 7735 -1912
rect 7706 -1919 7735 -1913
rect 8281 -1913 8287 -1912
rect 8304 -1898 8310 -1896
rect 8856 -1896 8885 -1890
rect 8856 -1898 8862 -1896
rect 8304 -1912 8316 -1898
rect 8850 -1912 8862 -1898
rect 8304 -1913 8310 -1912
rect 8281 -1919 8310 -1913
rect 8856 -1913 8862 -1912
rect 8879 -1898 8885 -1896
rect 9417 -1896 9446 -1890
rect 9417 -1898 9423 -1896
rect 8879 -1912 8891 -1898
rect 9411 -1912 9423 -1898
rect 8879 -1913 8885 -1912
rect 8856 -1919 8885 -1913
rect 9417 -1913 9423 -1912
rect 9440 -1898 9446 -1896
rect 9440 -1912 9452 -1898
rect 9440 -1913 9446 -1912
rect 9417 -1919 9446 -1913
rect -4549 -1964 240 -1950
rect -40 -2032 0 -2025
rect -40 -2058 -33 -2032
rect -7 -2038 0 -2032
rect 126 -2033 159 -2030
rect 126 -2038 130 -2033
rect -7 -2053 130 -2038
rect -7 -2058 0 -2053
rect -40 -2065 0 -2058
rect 126 -2059 130 -2053
rect 156 -2038 159 -2033
rect 156 -2052 228 -2038
rect 156 -2059 159 -2052
rect 126 -2062 159 -2059
rect 225 -2101 257 -2098
rect 225 -2127 228 -2101
rect 254 -2127 257 -2101
rect 225 -2130 257 -2127
rect 806 -2099 838 -2096
rect 806 -2125 809 -2099
rect 835 -2125 838 -2099
rect 806 -2128 838 -2125
rect 1378 -2100 1410 -2097
rect 1378 -2126 1381 -2100
rect 1407 -2126 1410 -2100
rect 1378 -2129 1410 -2126
rect 1956 -2102 1988 -2099
rect 1956 -2128 1959 -2102
rect 1985 -2128 1988 -2102
rect 1956 -2131 1988 -2128
rect 2531 -2102 2563 -2099
rect 2531 -2128 2534 -2102
rect 2560 -2128 2563 -2102
rect 2531 -2131 2563 -2128
rect 3102 -2104 3134 -2101
rect 3102 -2130 3105 -2104
rect 3131 -2130 3134 -2104
rect 3102 -2133 3134 -2130
rect 3679 -2103 3711 -2100
rect 3679 -2129 3682 -2103
rect 3708 -2129 3711 -2103
rect 3679 -2132 3711 -2129
rect 4259 -2102 4291 -2099
rect 4259 -2128 4262 -2102
rect 4288 -2128 4291 -2102
rect 4259 -2131 4291 -2128
rect 4829 -2101 4861 -2098
rect 4829 -2127 4832 -2101
rect 4858 -2127 4861 -2101
rect 4829 -2130 4861 -2127
rect 5406 -2103 5438 -2100
rect 5406 -2129 5409 -2103
rect 5435 -2129 5438 -2103
rect 5406 -2132 5438 -2129
rect 5980 -2101 6012 -2098
rect 5980 -2127 5983 -2101
rect 6009 -2127 6012 -2101
rect 5980 -2130 6012 -2127
rect 6553 -2102 6585 -2099
rect 6553 -2128 6556 -2102
rect 6582 -2128 6585 -2102
rect 6553 -2131 6585 -2128
rect 7130 -2103 7162 -2100
rect 7130 -2129 7133 -2103
rect 7159 -2129 7162 -2103
rect 7130 -2132 7162 -2129
rect 7706 -2103 7738 -2100
rect 7706 -2129 7709 -2103
rect 7735 -2129 7738 -2103
rect 7706 -2132 7738 -2129
rect 8279 -2105 8311 -2102
rect 8279 -2131 8282 -2105
rect 8308 -2131 8311 -2105
rect 8279 -2134 8311 -2131
rect 8854 -2105 8886 -2102
rect 8854 -2131 8857 -2105
rect 8883 -2131 8886 -2105
rect 8854 -2134 8886 -2131
rect 296 -2300 299 -2274
rect 325 -2280 328 -2274
rect 662 -2280 691 -2277
rect 749 -2280 752 -2274
rect 325 -2294 668 -2280
rect 325 -2300 328 -2294
rect 662 -2297 668 -2294
rect 685 -2294 752 -2280
rect 685 -2297 691 -2294
rect 662 -2300 691 -2297
rect 749 -2300 752 -2294
rect 778 -2300 781 -2274
rect 871 -2300 874 -2274
rect 900 -2280 903 -2274
rect 961 -2280 990 -2277
rect 1324 -2280 1327 -2274
rect 900 -2294 967 -2280
rect 900 -2300 903 -2294
rect 961 -2297 967 -2294
rect 984 -2294 1327 -2280
rect 984 -2297 990 -2294
rect 961 -2300 990 -2297
rect 1324 -2300 1327 -2294
rect 1353 -2300 1356 -2274
rect 1446 -2300 1449 -2274
rect 1475 -2280 1478 -2274
rect 1813 -2280 1842 -2277
rect 1899 -2280 1902 -2274
rect 1475 -2294 1819 -2280
rect 1475 -2300 1478 -2294
rect 1813 -2297 1819 -2294
rect 1836 -2294 1902 -2280
rect 1836 -2297 1842 -2294
rect 1813 -2300 1842 -2297
rect 1899 -2300 1902 -2294
rect 1928 -2300 1931 -2274
rect 2021 -2300 2024 -2274
rect 2050 -2280 2053 -2274
rect 2111 -2280 2140 -2277
rect 2474 -2280 2477 -2274
rect 2050 -2294 2117 -2280
rect 2050 -2300 2053 -2294
rect 2111 -2297 2117 -2294
rect 2134 -2294 2477 -2280
rect 2134 -2297 2140 -2294
rect 2111 -2300 2140 -2297
rect 2474 -2300 2477 -2294
rect 2503 -2300 2506 -2274
rect 2596 -2300 2599 -2274
rect 2625 -2280 2628 -2274
rect 2963 -2280 2992 -2277
rect 3049 -2280 3052 -2274
rect 2625 -2294 2969 -2280
rect 2625 -2300 2628 -2294
rect 2963 -2297 2969 -2294
rect 2986 -2294 3052 -2280
rect 2986 -2297 2992 -2294
rect 2963 -2300 2992 -2297
rect 3049 -2300 3052 -2294
rect 3078 -2300 3081 -2274
rect 3171 -2300 3174 -2274
rect 3200 -2280 3203 -2274
rect 3261 -2280 3290 -2277
rect 3624 -2280 3627 -2274
rect 3200 -2294 3267 -2280
rect 3200 -2300 3203 -2294
rect 3261 -2297 3267 -2294
rect 3284 -2294 3627 -2280
rect 3284 -2297 3290 -2294
rect 3261 -2300 3290 -2297
rect 3624 -2300 3627 -2294
rect 3653 -2300 3656 -2274
rect 3746 -2300 3749 -2274
rect 3775 -2280 3778 -2274
rect 4113 -2280 4142 -2277
rect 4199 -2280 4202 -2274
rect 3775 -2294 4119 -2280
rect 3775 -2300 3778 -2294
rect 4113 -2297 4119 -2294
rect 4136 -2294 4202 -2280
rect 4136 -2297 4142 -2294
rect 4113 -2300 4142 -2297
rect 4199 -2300 4202 -2294
rect 4228 -2300 4231 -2274
rect 4321 -2300 4324 -2274
rect 4350 -2280 4353 -2274
rect 4411 -2280 4440 -2277
rect 4774 -2280 4777 -2274
rect 4350 -2294 4417 -2280
rect 4350 -2300 4353 -2294
rect 4411 -2297 4417 -2294
rect 4434 -2294 4777 -2280
rect 4434 -2297 4440 -2294
rect 4411 -2300 4440 -2297
rect 4774 -2300 4777 -2294
rect 4803 -2300 4806 -2274
rect 4896 -2300 4899 -2274
rect 4925 -2280 4928 -2274
rect 5263 -2280 5292 -2277
rect 5349 -2280 5352 -2274
rect 4925 -2294 5269 -2280
rect 4925 -2300 4928 -2294
rect 5263 -2297 5269 -2294
rect 5286 -2294 5352 -2280
rect 5286 -2297 5292 -2294
rect 5263 -2300 5292 -2297
rect 5349 -2300 5352 -2294
rect 5378 -2300 5381 -2274
rect 5471 -2300 5474 -2274
rect 5500 -2280 5503 -2274
rect 5561 -2280 5590 -2277
rect 5924 -2280 5927 -2274
rect 5500 -2294 5567 -2280
rect 5500 -2300 5503 -2294
rect 5561 -2297 5567 -2294
rect 5584 -2294 5927 -2280
rect 5584 -2297 5590 -2294
rect 5561 -2300 5590 -2297
rect 5924 -2300 5927 -2294
rect 5953 -2300 5956 -2274
rect 6046 -2300 6049 -2274
rect 6075 -2280 6078 -2274
rect 6413 -2280 6442 -2277
rect 6499 -2280 6502 -2274
rect 6075 -2294 6419 -2280
rect 6075 -2300 6078 -2294
rect 6413 -2297 6419 -2294
rect 6436 -2294 6502 -2280
rect 6436 -2297 6442 -2294
rect 6413 -2300 6442 -2297
rect 6499 -2300 6502 -2294
rect 6528 -2300 6531 -2274
rect 6621 -2300 6624 -2274
rect 6650 -2280 6653 -2274
rect 6711 -2280 6740 -2277
rect 7074 -2280 7077 -2274
rect 6650 -2294 6717 -2280
rect 6650 -2300 6653 -2294
rect 6711 -2297 6717 -2294
rect 6734 -2294 7077 -2280
rect 6734 -2297 6740 -2294
rect 6711 -2300 6740 -2297
rect 7074 -2300 7077 -2294
rect 7103 -2300 7106 -2274
rect 7196 -2300 7199 -2274
rect 7225 -2280 7228 -2274
rect 7563 -2280 7592 -2277
rect 7649 -2280 7652 -2274
rect 7225 -2294 7569 -2280
rect 7225 -2300 7228 -2294
rect 7563 -2297 7569 -2294
rect 7586 -2294 7652 -2280
rect 7586 -2297 7592 -2294
rect 7563 -2300 7592 -2297
rect 7649 -2300 7652 -2294
rect 7678 -2300 7681 -2274
rect 7771 -2300 7774 -2274
rect 7800 -2280 7803 -2274
rect 7861 -2280 7890 -2277
rect 8224 -2280 8227 -2274
rect 7800 -2294 7867 -2280
rect 7800 -2300 7803 -2294
rect 7861 -2297 7867 -2294
rect 7884 -2294 8227 -2280
rect 7884 -2297 7890 -2294
rect 7861 -2300 7890 -2297
rect 8224 -2300 8227 -2294
rect 8253 -2300 8256 -2274
rect 8346 -2300 8349 -2274
rect 8375 -2280 8378 -2274
rect 8713 -2280 8742 -2277
rect 8799 -2280 8802 -2274
rect 8375 -2294 8719 -2280
rect 8375 -2300 8378 -2294
rect 8713 -2297 8719 -2294
rect 8736 -2294 8802 -2280
rect 8736 -2297 8742 -2294
rect 8713 -2300 8742 -2297
rect 8799 -2300 8802 -2294
rect 8828 -2300 8831 -2274
rect 8921 -2300 8924 -2274
rect 8950 -2280 8953 -2274
rect 9011 -2280 9040 -2277
rect 9374 -2280 9377 -2274
rect 8950 -2294 9017 -2280
rect 8950 -2300 8953 -2294
rect 9011 -2297 9017 -2294
rect 9034 -2294 9377 -2280
rect 9034 -2297 9040 -2294
rect 9011 -2300 9040 -2297
rect 9374 -2300 9377 -2294
rect 9403 -2300 9406 -2274
rect 806 -2322 846 -2315
rect 523 -2367 526 -2341
rect 552 -2367 555 -2341
rect 806 -2348 813 -2322
rect 839 -2348 846 -2322
rect 1955 -2323 1995 -2316
rect 806 -2355 846 -2348
rect 1098 -2368 1101 -2342
rect 1127 -2368 1130 -2342
rect 1673 -2373 1676 -2347
rect 1702 -2373 1705 -2347
rect 1955 -2349 1962 -2323
rect 1988 -2349 1995 -2323
rect 3098 -2324 3138 -2317
rect 1955 -2356 1995 -2349
rect 2248 -2373 2251 -2347
rect 2277 -2373 2280 -2347
rect 2823 -2373 2826 -2347
rect 2852 -2373 2855 -2347
rect 3098 -2350 3105 -2324
rect 3131 -2350 3138 -2324
rect 4255 -2325 4295 -2318
rect 3098 -2357 3138 -2350
rect 3398 -2373 3401 -2347
rect 3427 -2373 3430 -2347
rect 3973 -2373 3976 -2347
rect 4002 -2373 4005 -2347
rect 4255 -2351 4262 -2325
rect 4288 -2351 4295 -2325
rect 5395 -2323 5435 -2316
rect 4255 -2358 4295 -2351
rect 4548 -2373 4551 -2347
rect 4577 -2373 4580 -2347
rect 5123 -2373 5126 -2347
rect 5152 -2373 5155 -2347
rect 5395 -2349 5402 -2323
rect 5428 -2349 5435 -2323
rect 6563 -2323 6603 -2316
rect 5395 -2356 5435 -2349
rect 5698 -2373 5701 -2347
rect 5727 -2373 5730 -2347
rect 6273 -2373 6276 -2347
rect 6302 -2373 6305 -2347
rect 6563 -2349 6570 -2323
rect 6596 -2349 6603 -2323
rect 7708 -2323 7748 -2316
rect 6563 -2356 6603 -2349
rect 6848 -2373 6851 -2347
rect 6877 -2373 6880 -2347
rect 7423 -2373 7426 -2347
rect 7452 -2373 7455 -2347
rect 7708 -2349 7715 -2323
rect 7741 -2349 7748 -2323
rect 8865 -2321 8905 -2314
rect 8865 -2347 8872 -2321
rect 8898 -2347 8905 -2321
rect 7708 -2356 7748 -2349
rect 7998 -2373 8001 -2347
rect 8027 -2373 8030 -2347
rect 8573 -2373 8576 -2347
rect 8602 -2373 8605 -2347
rect 8865 -2354 8905 -2347
rect 9148 -2373 9151 -2347
rect 9177 -2373 9180 -2347
rect 730 -2421 770 -2414
rect 730 -2447 737 -2421
rect 763 -2447 770 -2421
rect 730 -2454 770 -2447
rect 885 -2421 925 -2414
rect 885 -2447 892 -2421
rect 918 -2447 925 -2421
rect 885 -2454 925 -2447
rect 1880 -2421 1920 -2414
rect 1880 -2447 1887 -2421
rect 1913 -2447 1920 -2421
rect 1880 -2454 1920 -2447
rect 2035 -2421 2075 -2414
rect 2035 -2447 2042 -2421
rect 2068 -2447 2075 -2421
rect 2035 -2454 2075 -2447
rect 3030 -2421 3070 -2414
rect 3030 -2447 3037 -2421
rect 3063 -2447 3070 -2421
rect 3030 -2454 3070 -2447
rect 3184 -2421 3224 -2414
rect 3184 -2447 3191 -2421
rect 3217 -2447 3224 -2421
rect 3184 -2454 3224 -2447
rect 4177 -2421 4217 -2414
rect 4177 -2447 4184 -2421
rect 4210 -2447 4217 -2421
rect 4177 -2454 4217 -2447
rect 4336 -2422 4376 -2415
rect 4336 -2448 4343 -2422
rect 4369 -2448 4376 -2422
rect -3927 -2484 -3924 -2458
rect -3898 -2461 -3895 -2458
rect 662 -2461 694 -2454
rect 4336 -2455 4376 -2448
rect 5329 -2421 5369 -2414
rect 5329 -2447 5336 -2421
rect 5362 -2447 5369 -2421
rect 5329 -2454 5369 -2447
rect 5484 -2421 5524 -2414
rect 5484 -2447 5491 -2421
rect 5517 -2447 5524 -2421
rect 5484 -2454 5524 -2447
rect 6480 -2422 6520 -2415
rect 6480 -2448 6487 -2422
rect 6513 -2448 6520 -2422
rect 6480 -2455 6520 -2448
rect 6633 -2422 6673 -2415
rect 6633 -2448 6640 -2422
rect 6666 -2448 6673 -2422
rect 6633 -2455 6673 -2448
rect 7631 -2421 7671 -2414
rect 7631 -2447 7638 -2421
rect 7664 -2447 7671 -2421
rect 7631 -2454 7671 -2447
rect 7784 -2421 7824 -2414
rect 7784 -2447 7791 -2421
rect 7817 -2447 7824 -2421
rect 7784 -2454 7824 -2447
rect 8780 -2420 8820 -2414
rect 8780 -2446 8787 -2420
rect 8813 -2446 8820 -2420
rect 8780 -2454 8820 -2446
rect 8932 -2421 8972 -2413
rect 8932 -2447 8939 -2421
rect 8965 -2447 8972 -2421
rect 8932 -2454 8972 -2447
rect -3898 -2462 694 -2461
rect -3898 -2475 669 -2462
rect -3898 -2484 -3895 -2475
rect 662 -2479 669 -2475
rect 686 -2479 694 -2462
rect 662 -2485 694 -2479
rect 1154 -2491 1194 -2484
rect 461 -2498 501 -2491
rect 461 -2524 468 -2498
rect 494 -2524 501 -2498
rect 1154 -2517 1161 -2491
rect 1187 -2517 1194 -2491
rect 1154 -2524 1194 -2517
rect 1610 -2490 1650 -2483
rect 1610 -2516 1617 -2490
rect 1643 -2516 1650 -2490
rect 1610 -2523 1650 -2516
rect 2303 -2495 2343 -2488
rect 2303 -2521 2310 -2495
rect 2336 -2521 2343 -2495
rect 461 -2531 501 -2524
rect 2303 -2528 2343 -2521
rect 2762 -2496 2802 -2489
rect 2762 -2522 2769 -2496
rect 2795 -2522 2802 -2496
rect 2762 -2529 2802 -2522
rect 3454 -2494 3494 -2487
rect 3454 -2520 3461 -2494
rect 3487 -2520 3494 -2494
rect 3454 -2527 3494 -2520
rect 3912 -2496 3952 -2489
rect 3912 -2522 3919 -2496
rect 3945 -2522 3952 -2496
rect 3912 -2529 3952 -2522
rect 4603 -2498 4643 -2491
rect 4603 -2524 4610 -2498
rect 4636 -2524 4643 -2498
rect 4603 -2531 4643 -2524
rect 5061 -2492 5101 -2485
rect 5061 -2518 5068 -2492
rect 5094 -2518 5101 -2492
rect 5061 -2525 5101 -2518
rect 5754 -2494 5794 -2487
rect 5754 -2520 5761 -2494
rect 5787 -2520 5794 -2494
rect 5754 -2527 5794 -2520
rect 6211 -2490 6251 -2483
rect 6211 -2516 6218 -2490
rect 6244 -2516 6251 -2490
rect 6211 -2523 6251 -2516
rect 6903 -2494 6943 -2487
rect 6903 -2520 6910 -2494
rect 6936 -2520 6943 -2494
rect 6903 -2527 6943 -2520
rect 7361 -2494 7401 -2487
rect 7361 -2520 7368 -2494
rect 7394 -2520 7401 -2494
rect 7361 -2527 7401 -2520
rect 8053 -2497 8093 -2490
rect 8053 -2523 8060 -2497
rect 8086 -2523 8093 -2497
rect 8053 -2530 8093 -2523
rect 8511 -2495 8551 -2489
rect 8511 -2521 8518 -2495
rect 8544 -2521 8551 -2495
rect 8511 -2529 8551 -2521
rect 9203 -2491 9239 -2487
rect 9203 -2521 9206 -2491
rect 9236 -2521 9239 -2491
rect 9203 -2525 9239 -2521
rect -2747 -2566 -2744 -2540
rect -2718 -2545 -2715 -2540
rect 963 -2545 991 -2540
rect -2718 -2546 991 -2545
rect -2718 -2562 968 -2546
rect -2718 -2566 -2715 -2562
rect 963 -2563 968 -2562
rect 985 -2563 991 -2546
rect 9012 -2542 9041 -2540
rect 13529 -2542 13532 -2537
rect 9012 -2543 13532 -2542
rect 9012 -2560 9018 -2543
rect 9035 -2559 13532 -2543
rect 9035 -2560 9041 -2559
rect 9012 -2563 9041 -2560
rect 13529 -2563 13532 -2559
rect 13558 -2563 13561 -2537
rect 963 -2569 991 -2563
rect 12586 -2587 12612 -2584
rect 8712 -2592 8741 -2590
rect 8712 -2593 12586 -2592
rect -1568 -2629 -1565 -2603
rect -1539 -2608 -1536 -2603
rect 1812 -2608 1841 -2602
rect -1539 -2609 1841 -2608
rect -1539 -2625 1818 -2609
rect -1539 -2629 -1536 -2625
rect 1812 -2626 1818 -2625
rect 1835 -2626 1841 -2609
rect 8712 -2610 8718 -2593
rect 8735 -2609 12586 -2593
rect 8735 -2610 8741 -2609
rect 8712 -2613 8741 -2610
rect 12586 -2616 12612 -2613
rect 1812 -2631 1841 -2626
rect 11423 -2637 11449 -2634
rect 7862 -2642 7891 -2640
rect 7862 -2643 11423 -2642
rect 7862 -2660 7868 -2643
rect 7885 -2659 11423 -2643
rect 7885 -2660 7891 -2659
rect 7862 -2663 7891 -2660
rect 11423 -2666 11449 -2663
rect -390 -2704 -387 -2678
rect -361 -2683 -358 -2678
rect 2112 -2683 2141 -2681
rect -361 -2684 2141 -2683
rect -361 -2700 2118 -2684
rect -361 -2704 -358 -2700
rect 2112 -2701 2118 -2700
rect 2135 -2701 2141 -2684
rect 2112 -2704 2141 -2701
rect 10210 -2700 10236 -2697
rect 7562 -2705 7591 -2703
rect 7562 -2706 10210 -2705
rect 7562 -2723 7568 -2706
rect 7585 -2722 10210 -2706
rect 7585 -2723 7591 -2722
rect 7562 -2726 7591 -2723
rect 10210 -2729 10236 -2726
rect 808 -2775 811 -2749
rect 837 -2754 840 -2749
rect 2962 -2754 2991 -2752
rect 837 -2755 2991 -2754
rect 837 -2771 2968 -2755
rect 837 -2775 840 -2771
rect 2962 -2772 2968 -2771
rect 2985 -2772 2991 -2755
rect 9036 -2763 9062 -2760
rect 2962 -2775 2991 -2772
rect 6715 -2768 6738 -2763
rect 6715 -2769 9036 -2768
rect 6715 -2786 6718 -2769
rect 6735 -2785 9036 -2769
rect 6735 -2786 6738 -2785
rect 6715 -2792 6738 -2786
rect 9036 -2792 9062 -2789
rect 1975 -2855 1978 -2829
rect 2004 -2834 2007 -2829
rect 3262 -2834 3291 -2832
rect 2004 -2835 3291 -2834
rect 2004 -2851 3268 -2835
rect 2004 -2855 2007 -2851
rect 3262 -2852 3268 -2851
rect 3285 -2852 3291 -2835
rect 3262 -2855 3291 -2852
rect 6412 -2840 6441 -2838
rect 7845 -2840 7848 -2835
rect 6412 -2841 7848 -2840
rect 6412 -2858 6418 -2841
rect 6435 -2857 7848 -2841
rect 6435 -2858 6441 -2857
rect 6412 -2861 6441 -2858
rect 7845 -2861 7848 -2857
rect 7874 -2861 7877 -2835
rect 3137 -2913 3163 -2910
rect 4112 -2918 4141 -2916
rect 3163 -2919 4141 -2918
rect 3163 -2935 4118 -2919
rect 4112 -2936 4118 -2935
rect 4135 -2936 4141 -2919
rect 4112 -2939 4141 -2936
rect 5562 -2920 5591 -2918
rect 6643 -2920 6646 -2915
rect 5562 -2921 6646 -2920
rect 5562 -2938 5568 -2921
rect 5585 -2937 6646 -2921
rect 5585 -2938 5591 -2937
rect 3137 -2942 3163 -2939
rect 5562 -2941 5591 -2938
rect 6643 -2941 6646 -2937
rect 6672 -2941 6675 -2915
rect 4308 -3010 4311 -2984
rect 4337 -2989 4340 -2984
rect 4412 -2989 4441 -2987
rect 4337 -2990 4441 -2989
rect 4337 -3006 4418 -2990
rect 4337 -3010 4340 -3006
rect 4412 -3007 4418 -3006
rect 4435 -3007 4441 -2990
rect 4412 -3010 4441 -3007
rect 5262 -3007 5291 -3005
rect 5493 -3007 5496 -3002
rect 5262 -3008 5496 -3007
rect 5262 -3025 5268 -3008
rect 5285 -3024 5496 -3008
rect 5285 -3025 5291 -3024
rect 5262 -3028 5291 -3025
rect 5493 -3028 5496 -3024
rect 5522 -3028 5525 -3002
rect -3991 -3151 -3988 -3125
rect -3962 -3131 -3959 -3125
rect -3962 -3145 -3830 -3131
rect -3196 -3145 -2694 -3131
rect -2049 -3145 -1512 -3131
rect -864 -3145 -330 -3131
rect 317 -3145 850 -3131
rect 1498 -3145 2032 -3131
rect 2680 -3145 3214 -3131
rect 3862 -3145 4396 -3131
rect 5043 -3145 5578 -3131
rect 6223 -3145 6760 -3131
rect 7408 -3145 7942 -3131
rect 8590 -3145 9126 -3131
rect 9774 -3145 10310 -3131
rect 10958 -3145 11497 -3131
rect 12145 -3145 12684 -3131
rect 13332 -3145 13585 -3131
rect -3962 -3151 -3959 -3145
rect -3660 -3589 -3631 -3583
rect -3660 -3606 -3654 -3589
rect -3637 -3590 -3631 -3589
rect -3151 -3590 -3148 -3584
rect -3637 -3604 -3148 -3590
rect -3637 -3606 -3631 -3604
rect -3660 -3612 -3631 -3606
rect -3151 -3610 -3148 -3604
rect -3122 -3610 -3119 -3584
rect -2487 -3589 -2458 -3583
rect -2487 -3606 -2481 -3589
rect -2464 -3590 -2458 -3589
rect -1996 -3590 -1993 -3584
rect -2464 -3604 -1993 -3590
rect -2464 -3606 -2458 -3604
rect -2487 -3612 -2458 -3606
rect -1996 -3610 -1993 -3604
rect -1967 -3610 -1964 -3584
rect -1312 -3589 -1289 -3583
rect -1312 -3606 -1309 -3589
rect -1292 -3590 -1289 -3589
rect -827 -3590 -824 -3584
rect -1292 -3604 -824 -3590
rect -1292 -3606 -1289 -3604
rect -1312 -3612 -1289 -3606
rect -827 -3610 -824 -3604
rect -798 -3610 -795 -3584
rect -134 -3589 -105 -3583
rect -134 -3606 -128 -3589
rect -111 -3590 -105 -3589
rect 364 -3590 367 -3584
rect -111 -3604 367 -3590
rect -111 -3606 -105 -3604
rect -134 -3612 -105 -3606
rect 364 -3610 367 -3604
rect 393 -3610 396 -3584
rect 1052 -3589 1081 -3583
rect 1052 -3606 1058 -3589
rect 1075 -3590 1081 -3589
rect 1541 -3590 1544 -3584
rect 1075 -3604 1544 -3590
rect 1075 -3606 1081 -3604
rect 1052 -3612 1081 -3606
rect 1541 -3610 1544 -3604
rect 1570 -3610 1573 -3584
rect 2236 -3589 2265 -3583
rect 2236 -3606 2242 -3589
rect 2259 -3590 2265 -3589
rect 2718 -3590 2721 -3584
rect 2259 -3604 2721 -3590
rect 2259 -3606 2265 -3604
rect 2236 -3612 2265 -3606
rect 2718 -3610 2721 -3604
rect 2747 -3610 2750 -3584
rect 3404 -3589 3433 -3583
rect 3404 -3606 3410 -3589
rect 3427 -3590 3433 -3589
rect 3900 -3590 3903 -3584
rect 3427 -3604 3903 -3590
rect 3427 -3606 3433 -3604
rect 3404 -3612 3433 -3606
rect 3900 -3610 3903 -3604
rect 3929 -3610 3932 -3584
rect 4593 -3589 4622 -3583
rect 4593 -3606 4599 -3589
rect 4616 -3590 4622 -3589
rect 5086 -3590 5089 -3584
rect 4616 -3604 5089 -3590
rect 4616 -3606 4622 -3604
rect 4593 -3612 4622 -3606
rect 5086 -3610 5089 -3604
rect 5115 -3610 5118 -3584
rect 5771 -3589 5800 -3583
rect 5771 -3606 5777 -3589
rect 5794 -3590 5800 -3589
rect 6265 -3590 6268 -3584
rect 5794 -3604 6268 -3590
rect 5794 -3606 5800 -3604
rect 5771 -3612 5800 -3606
rect 6265 -3610 6268 -3604
rect 6294 -3610 6297 -3584
rect 6960 -3589 6989 -3583
rect 6960 -3606 6966 -3589
rect 6983 -3590 6989 -3589
rect 7453 -3590 7456 -3584
rect 6983 -3604 7456 -3590
rect 6983 -3606 6989 -3604
rect 6960 -3612 6989 -3606
rect 7453 -3610 7456 -3604
rect 7482 -3610 7485 -3584
rect 8126 -3589 8155 -3583
rect 8126 -3606 8132 -3589
rect 8149 -3590 8155 -3589
rect 8626 -3590 8629 -3584
rect 8149 -3604 8629 -3590
rect 8149 -3606 8155 -3604
rect 8126 -3612 8155 -3606
rect 8626 -3610 8629 -3604
rect 8655 -3610 8658 -3584
rect 9328 -3589 9357 -3583
rect 9328 -3606 9334 -3589
rect 9351 -3590 9357 -3589
rect 9808 -3590 9811 -3584
rect 9351 -3604 9811 -3590
rect 9351 -3606 9357 -3604
rect 9328 -3612 9357 -3606
rect 9808 -3610 9811 -3604
rect 9837 -3610 9840 -3584
rect 10501 -3589 10530 -3583
rect 10501 -3606 10507 -3589
rect 10524 -3590 10530 -3589
rect 10997 -3590 11000 -3584
rect 10524 -3604 11000 -3590
rect 10524 -3606 10530 -3604
rect 10501 -3612 10530 -3606
rect 10997 -3610 11000 -3604
rect 11026 -3610 11029 -3584
rect 11673 -3589 11702 -3583
rect 11673 -3606 11679 -3589
rect 11696 -3590 11702 -3589
rect 12192 -3590 12195 -3584
rect 11696 -3604 12195 -3590
rect 11696 -3606 11702 -3604
rect 11673 -3612 11702 -3606
rect 12192 -3610 12195 -3604
rect 12221 -3610 12224 -3584
rect 12889 -3589 12918 -3583
rect 12889 -3606 12895 -3589
rect 12912 -3590 12918 -3589
rect 13368 -3590 13371 -3584
rect 12912 -3604 13371 -3590
rect 12912 -3606 12918 -3604
rect 12889 -3612 12918 -3606
rect 13368 -3610 13371 -3604
rect 13397 -3610 13400 -3584
rect 13791 -3589 13820 -3583
rect 13791 -3606 13797 -3589
rect 13814 -3590 13820 -3589
rect 14272 -3590 14275 -3584
rect 13814 -3604 14275 -3590
rect 13814 -3606 13820 -3604
rect 13791 -3612 13820 -3606
rect 14272 -3610 14275 -3604
rect 14301 -3610 14304 -3584
rect -4057 -3654 -4054 -3628
rect -4028 -3634 -4025 -3628
rect -4028 -3648 -3829 -3634
rect -3196 -3648 -2694 -3634
rect -2046 -3648 -1512 -3634
rect -864 -3648 -331 -3634
rect 317 -3648 850 -3634
rect 1498 -3648 2032 -3634
rect 2680 -3648 3214 -3634
rect 3861 -3648 4397 -3634
rect 5044 -3648 5578 -3634
rect 6226 -3648 6760 -3634
rect 7407 -3648 7942 -3634
rect 8590 -3648 9126 -3634
rect 9774 -3648 10310 -3634
rect 10955 -3648 11497 -3634
rect 12145 -3648 12684 -3634
rect 13332 -3648 13585 -3634
rect -4028 -3654 -4025 -3648
rect -4123 -3694 -4120 -3668
rect -4094 -3674 -4091 -3668
rect -4094 -3688 -3830 -3674
rect -3196 -3688 -2694 -3674
rect -2046 -3688 -1512 -3674
rect -865 -3688 -331 -3674
rect 313 -3688 850 -3674
rect 1498 -3688 2032 -3674
rect 2680 -3688 3214 -3674
rect 3862 -3688 4396 -3674
rect 5042 -3688 5578 -3674
rect 6226 -3688 6760 -3674
rect 7406 -3688 7942 -3674
rect 8590 -3688 9126 -3674
rect 9770 -3688 10310 -3674
rect 10954 -3688 11497 -3674
rect 12141 -3688 12684 -3674
rect 13330 -3688 13585 -3674
rect -4094 -3694 -4091 -3688
rect -3930 -4131 -3892 -4128
rect -3930 -4163 -3927 -4131
rect -3895 -4140 -3892 -4131
rect -2743 -4135 -2717 -4132
rect -3895 -4154 -3844 -4140
rect -3895 -4163 -3892 -4154
rect -3930 -4166 -3892 -4163
rect -2717 -4156 -2694 -4139
rect -1567 -4161 -1564 -4135
rect -1538 -4139 -1535 -4135
rect -1538 -4156 -1512 -4139
rect -1538 -4161 -1535 -4156
rect -389 -4161 -386 -4135
rect -360 -4139 -357 -4135
rect -360 -4156 -331 -4139
rect -360 -4161 -357 -4156
rect 809 -4161 812 -4135
rect 838 -4139 841 -4135
rect 838 -4154 850 -4139
rect 838 -4161 841 -4154
rect 1976 -4160 1979 -4134
rect 2005 -4138 2008 -4134
rect 2005 -4155 2032 -4138
rect 2005 -4160 2008 -4155
rect 3135 -4159 3138 -4133
rect 3164 -4137 3167 -4133
rect 3164 -4154 3214 -4137
rect 3164 -4159 3167 -4154
rect 4309 -4159 4312 -4133
rect 4338 -4137 4341 -4133
rect 4338 -4154 4396 -4137
rect 4338 -4159 4341 -4154
rect 5494 -4159 5497 -4133
rect 5523 -4137 5526 -4133
rect 9037 -4135 9063 -4132
rect 13533 -4134 13559 -4131
rect 5523 -4154 5578 -4137
rect 5523 -4159 5526 -4154
rect 6644 -4161 6647 -4135
rect 6673 -4139 6676 -4135
rect 6673 -4156 6760 -4139
rect 6673 -4161 6676 -4156
rect 7846 -4161 7849 -4135
rect 7875 -4139 7878 -4135
rect 7875 -4156 7942 -4139
rect 7875 -4161 7878 -4156
rect 9063 -4156 9126 -4139
rect 10208 -4161 10211 -4135
rect 10237 -4139 10240 -4135
rect 10237 -4156 10310 -4139
rect 10237 -4161 10240 -4156
rect 11421 -4160 11424 -4134
rect 11450 -4138 11453 -4134
rect 11450 -4155 11497 -4138
rect 11450 -4160 11453 -4155
rect 12584 -4161 12587 -4135
rect 12613 -4139 12616 -4135
rect 12613 -4156 12684 -4139
rect 12613 -4161 12616 -4156
rect 13559 -4155 13585 -4138
rect -2743 -4164 -2717 -4161
rect 9037 -4164 9063 -4161
rect 13533 -4163 13559 -4160
rect -4181 -4372 -4178 -4346
rect -4152 -4352 -4149 -4346
rect -3916 -4352 -3913 -4346
rect -4152 -4366 -3913 -4352
rect -4152 -4372 -4149 -4366
rect -3916 -4372 -3913 -4366
rect -3887 -4352 -3884 -4346
rect -3887 -4366 -3830 -4352
rect -3218 -4366 13585 -4352
rect -3887 -4372 -3884 -4366
rect -3221 -4450 -3192 -4448
rect -2071 -4450 -2042 -4447
rect -889 -4450 -860 -4447
rect 292 -4450 321 -4447
rect 1473 -4450 1502 -4447
rect 2655 -4450 2684 -4447
rect 3837 -4450 3866 -4447
rect 5019 -4450 5048 -4447
rect 6201 -4450 6230 -4447
rect 7383 -4450 7412 -4447
rect 8565 -4450 8594 -4447
rect 9749 -4450 9778 -4447
rect 10933 -4450 10962 -4447
rect 12120 -4450 12149 -4447
rect 13307 -4450 13336 -4447
rect 14211 -4450 14234 -4444
rect 14443 -4450 14446 -4445
rect -3221 -4451 -2065 -4450
rect -3221 -4468 -3215 -4451
rect -3198 -4467 -2065 -4451
rect -2048 -4467 -883 -4450
rect -866 -4467 298 -4450
rect 315 -4467 1479 -4450
rect 1496 -4467 2661 -4450
rect 2678 -4467 3843 -4450
rect 3860 -4467 5025 -4450
rect 5042 -4467 6207 -4450
rect 6224 -4467 7389 -4450
rect 7406 -4467 8571 -4450
rect 8588 -4467 9755 -4450
rect 9772 -4467 10939 -4450
rect 10956 -4467 12126 -4450
rect 12143 -4467 13313 -4450
rect 13330 -4467 14214 -4450
rect 14231 -4467 14446 -4450
rect -3198 -4468 -3192 -4467
rect -3221 -4471 -3192 -4468
rect -2071 -4470 -2042 -4467
rect -889 -4470 -860 -4467
rect 292 -4470 321 -4467
rect 1473 -4470 1502 -4467
rect 2655 -4470 2684 -4467
rect 3837 -4470 3866 -4467
rect 5019 -4470 5048 -4467
rect 6201 -4470 6230 -4467
rect 7383 -4470 7412 -4467
rect 8565 -4470 8594 -4467
rect 9749 -4470 9778 -4467
rect 10933 -4470 10962 -4467
rect 12120 -4470 12149 -4467
rect 13307 -4470 13336 -4467
rect 14211 -4473 14234 -4467
rect 14443 -4471 14446 -4467
rect 14472 -4471 14475 -4445
rect -3221 -4539 -3192 -4537
rect -2071 -4539 -2042 -4536
rect 292 -4539 321 -4536
rect 1473 -4539 1502 -4536
rect 2655 -4539 2684 -4536
rect 3837 -4539 3866 -4536
rect 5019 -4539 5048 -4536
rect 6201 -4539 6230 -4536
rect 7383 -4539 7412 -4536
rect 8565 -4539 8594 -4536
rect 9749 -4539 9778 -4536
rect 10933 -4539 10962 -4537
rect 12120 -4539 12149 -4536
rect 13307 -4539 13336 -4536
rect 14208 -4539 14237 -4536
rect 14499 -4539 14502 -4534
rect -3221 -4540 -2065 -4539
rect -3221 -4557 -3215 -4540
rect -3198 -4556 -2065 -4540
rect -2048 -4542 298 -4539
rect -2048 -4556 -883 -4542
rect -3198 -4557 -3192 -4556
rect -3221 -4560 -3192 -4557
rect -2071 -4559 -2042 -4556
rect -889 -4559 -883 -4556
rect -866 -4556 298 -4542
rect 315 -4556 1479 -4539
rect 1496 -4556 2661 -4539
rect 2678 -4556 3843 -4539
rect 3860 -4556 5025 -4539
rect 5042 -4556 6207 -4539
rect 6224 -4556 7389 -4539
rect 7406 -4556 8571 -4539
rect 8588 -4556 9755 -4539
rect 9772 -4540 12126 -4539
rect 9772 -4556 10939 -4540
rect -866 -4559 -860 -4556
rect 292 -4559 321 -4556
rect 1473 -4559 1502 -4556
rect 2655 -4559 2684 -4556
rect 3837 -4559 3866 -4556
rect 5019 -4559 5048 -4556
rect 6201 -4559 6230 -4556
rect 7383 -4559 7412 -4556
rect 8565 -4559 8594 -4556
rect 9749 -4559 9778 -4556
rect 10933 -4557 10939 -4556
rect 10956 -4556 12126 -4540
rect 12143 -4556 13313 -4539
rect 13330 -4556 14214 -4539
rect 14231 -4556 14502 -4539
rect 10956 -4557 10962 -4556
rect -889 -4562 -860 -4559
rect 10933 -4560 10962 -4557
rect 12120 -4559 12149 -4556
rect 13307 -4559 13336 -4556
rect 14208 -4559 14237 -4556
rect 14499 -4560 14502 -4556
rect 14528 -4560 14531 -4534
rect -3916 -4662 -3913 -4636
rect -3887 -4642 -3884 -4636
rect -3887 -4656 -3824 -4642
rect -3196 -4656 -2694 -4642
rect -2046 -4656 -1512 -4642
rect -864 -4656 -331 -4642
rect 317 -4656 850 -4642
rect 1498 -4656 2032 -4642
rect 2680 -4656 3214 -4642
rect 3862 -4656 4396 -4642
rect 5044 -4656 5578 -4642
rect 6226 -4656 6760 -4642
rect 7408 -4656 7942 -4642
rect 8590 -4656 9126 -4642
rect 9774 -4656 10310 -4642
rect 10958 -4656 11497 -4642
rect 12145 -4656 12684 -4642
rect 13332 -4656 13585 -4642
rect -3887 -4662 -3884 -4656
rect -4123 -5340 -4120 -5314
rect -4094 -5320 -4091 -5314
rect -4094 -5334 -3828 -5320
rect -3197 -5334 -2694 -5320
rect -2047 -5334 -1512 -5320
rect -864 -5334 -331 -5320
rect 317 -5334 850 -5320
rect 1498 -5334 2032 -5320
rect 2670 -5334 3214 -5320
rect 3859 -5334 4396 -5320
rect 5044 -5334 5578 -5320
rect 6226 -5334 6760 -5320
rect 7408 -5334 7942 -5320
rect 8588 -5334 9126 -5320
rect 9772 -5334 10310 -5320
rect 10954 -5334 11499 -5320
rect 12141 -5334 12684 -5320
rect 13332 -5334 13585 -5320
rect -4094 -5340 -4091 -5334
rect -4057 -5380 -4054 -5354
rect -4028 -5360 -4025 -5354
rect -4028 -5374 -3830 -5360
rect -3196 -5374 -2692 -5360
rect -2046 -5374 -1512 -5360
rect -864 -5374 -330 -5360
rect 317 -5374 850 -5360
rect 1498 -5374 2032 -5360
rect 2680 -5374 3214 -5360
rect 3862 -5374 4396 -5360
rect 5044 -5374 5578 -5360
rect 6226 -5374 6760 -5360
rect 7408 -5374 7942 -5360
rect 8590 -5374 9126 -5360
rect 9774 -5374 10310 -5360
rect 10958 -5374 11497 -5360
rect 12145 -5374 12684 -5360
rect 13332 -5374 13585 -5360
rect -4028 -5380 -4025 -5374
rect -3638 -5401 -3609 -5398
rect -3638 -5418 -3632 -5401
rect -3615 -5403 -3609 -5401
rect -3110 -5403 -3107 -5397
rect -3615 -5417 -3107 -5403
rect -3615 -5418 -3609 -5417
rect -3638 -5421 -3609 -5418
rect -3110 -5423 -3107 -5417
rect -3081 -5423 -3078 -5397
rect -2507 -5402 -2478 -5396
rect -2507 -5419 -2501 -5402
rect -2484 -5403 -2478 -5402
rect -1956 -5403 -1953 -5397
rect -2484 -5417 -1953 -5403
rect -2484 -5419 -2478 -5417
rect -2507 -5425 -2478 -5419
rect -1956 -5423 -1953 -5417
rect -1927 -5423 -1924 -5397
rect -1326 -5402 -1297 -5396
rect -1326 -5419 -1320 -5402
rect -1303 -5403 -1297 -5402
rect -787 -5403 -784 -5397
rect -1303 -5417 -784 -5403
rect -1303 -5419 -1297 -5417
rect -1326 -5425 -1297 -5419
rect -787 -5423 -784 -5417
rect -758 -5423 -755 -5397
rect -154 -5402 -125 -5396
rect -154 -5419 -148 -5402
rect -131 -5403 -125 -5402
rect 404 -5403 407 -5397
rect -131 -5417 407 -5403
rect -131 -5419 -125 -5417
rect -154 -5425 -125 -5419
rect 404 -5423 407 -5417
rect 433 -5423 436 -5397
rect 1024 -5402 1053 -5396
rect 1024 -5419 1030 -5402
rect 1047 -5403 1053 -5402
rect 1581 -5403 1584 -5397
rect 1047 -5417 1584 -5403
rect 1047 -5419 1053 -5417
rect 1024 -5425 1053 -5419
rect 1581 -5423 1584 -5417
rect 1610 -5423 1613 -5397
rect 2212 -5402 2241 -5396
rect 2212 -5419 2218 -5402
rect 2235 -5403 2241 -5402
rect 2758 -5403 2761 -5397
rect 2235 -5417 2761 -5403
rect 2235 -5419 2241 -5417
rect 2212 -5425 2241 -5419
rect 2758 -5423 2761 -5417
rect 2787 -5423 2790 -5397
rect 3403 -5402 3432 -5396
rect 3403 -5419 3409 -5402
rect 3426 -5403 3432 -5402
rect 3940 -5403 3943 -5397
rect 3426 -5417 3943 -5403
rect 3426 -5419 3432 -5417
rect 3403 -5425 3432 -5419
rect 3940 -5423 3943 -5417
rect 3969 -5423 3972 -5397
rect 4588 -5402 4611 -5396
rect 4588 -5419 4591 -5402
rect 4608 -5403 4611 -5402
rect 5126 -5403 5129 -5397
rect 4608 -5417 5129 -5403
rect 4608 -5419 4611 -5417
rect 4588 -5425 4611 -5419
rect 5126 -5423 5129 -5417
rect 5155 -5423 5158 -5397
rect 5754 -5402 5783 -5396
rect 5754 -5419 5760 -5402
rect 5777 -5403 5783 -5402
rect 6305 -5403 6308 -5397
rect 5777 -5417 6308 -5403
rect 5777 -5419 5783 -5417
rect 5754 -5425 5783 -5419
rect 6305 -5423 6308 -5417
rect 6334 -5423 6337 -5397
rect 6942 -5402 6971 -5396
rect 6942 -5419 6948 -5402
rect 6965 -5403 6971 -5402
rect 7493 -5403 7496 -5397
rect 6965 -5417 7496 -5403
rect 6965 -5419 6971 -5417
rect 6942 -5425 6971 -5419
rect 7493 -5423 7496 -5417
rect 7522 -5423 7525 -5397
rect 8121 -5402 8150 -5396
rect 8121 -5419 8127 -5402
rect 8144 -5403 8150 -5402
rect 8666 -5403 8669 -5397
rect 8144 -5417 8669 -5403
rect 8144 -5419 8150 -5417
rect 8121 -5425 8150 -5419
rect 8666 -5423 8669 -5417
rect 8695 -5423 8698 -5397
rect 9309 -5402 9338 -5396
rect 9309 -5419 9315 -5402
rect 9332 -5403 9338 -5402
rect 9848 -5403 9851 -5397
rect 9332 -5417 9851 -5403
rect 9332 -5419 9338 -5417
rect 9309 -5425 9338 -5419
rect 9848 -5423 9851 -5417
rect 9877 -5423 9880 -5397
rect 10486 -5402 10515 -5396
rect 10486 -5419 10492 -5402
rect 10509 -5403 10515 -5402
rect 11037 -5403 11040 -5397
rect 10509 -5417 11040 -5403
rect 10509 -5419 10515 -5417
rect 10486 -5425 10515 -5419
rect 11037 -5423 11040 -5417
rect 11066 -5423 11069 -5397
rect 11664 -5402 11693 -5396
rect 11664 -5419 11670 -5402
rect 11687 -5403 11693 -5402
rect 12232 -5403 12235 -5397
rect 11687 -5417 12235 -5403
rect 11687 -5419 11693 -5417
rect 11664 -5425 11693 -5419
rect 12232 -5423 12235 -5417
rect 12261 -5423 12264 -5397
rect 12845 -5402 12874 -5396
rect 12845 -5419 12851 -5402
rect 12868 -5403 12874 -5402
rect 13408 -5403 13411 -5397
rect 12868 -5417 13411 -5403
rect 12868 -5419 12874 -5417
rect 12845 -5425 12874 -5419
rect 13408 -5423 13411 -5417
rect 13437 -5423 13440 -5397
rect 13772 -5402 13801 -5396
rect 13772 -5419 13778 -5402
rect 13795 -5403 13801 -5402
rect 14312 -5403 14315 -5397
rect 13795 -5417 14315 -5403
rect 13795 -5419 13801 -5417
rect 13772 -5425 13801 -5419
rect 14312 -5423 14315 -5417
rect 14341 -5423 14344 -5397
rect -3990 -5883 -3987 -5857
rect -3961 -5863 -3958 -5857
rect -3961 -5878 -3829 -5863
rect -3197 -5878 -2694 -5863
rect -2047 -5878 -1512 -5863
rect -865 -5878 -331 -5863
rect 316 -5878 850 -5863
rect 1497 -5878 2032 -5863
rect 2677 -5878 3214 -5863
rect 3861 -5878 4396 -5863
rect 5042 -5878 5578 -5863
rect 6225 -5878 6760 -5863
rect 7406 -5878 7942 -5863
rect 8584 -5878 9126 -5863
rect 9773 -5878 10311 -5863
rect 10956 -5878 11497 -5863
rect 12144 -5878 12684 -5863
rect 13331 -5878 13585 -5863
rect -3961 -5883 -3958 -5878
rect -3637 -6322 -3614 -6316
rect -3637 -6339 -3634 -6322
rect -3617 -6323 -3614 -6322
rect -3070 -6323 -3067 -6317
rect -3617 -6337 -3067 -6323
rect -3617 -6339 -3614 -6337
rect -3637 -6345 -3614 -6339
rect -3070 -6343 -3067 -6337
rect -3041 -6343 -3038 -6317
rect -2493 -6322 -2463 -6316
rect -2493 -6339 -2486 -6322
rect -2469 -6323 -2463 -6322
rect -1914 -6323 -1911 -6317
rect -2469 -6337 -1911 -6323
rect -2469 -6339 -2463 -6337
rect -2493 -6345 -2463 -6339
rect -1914 -6343 -1911 -6337
rect -1885 -6343 -1882 -6317
rect -1311 -6322 -1282 -6316
rect -1311 -6339 -1305 -6322
rect -1288 -6323 -1282 -6322
rect -745 -6323 -742 -6317
rect -1288 -6337 -742 -6323
rect -1288 -6339 -1282 -6337
rect -1311 -6345 -1282 -6339
rect -745 -6343 -742 -6337
rect -716 -6343 -713 -6317
rect -136 -6322 -107 -6316
rect -136 -6339 -130 -6322
rect -113 -6323 -107 -6322
rect 446 -6323 449 -6317
rect -113 -6337 449 -6323
rect -113 -6339 -107 -6337
rect -136 -6344 -107 -6339
rect 446 -6343 449 -6337
rect 475 -6343 478 -6317
rect 1052 -6322 1081 -6316
rect 1052 -6339 1058 -6322
rect 1075 -6323 1081 -6322
rect 1623 -6323 1626 -6317
rect 1075 -6337 1626 -6323
rect 1075 -6339 1081 -6337
rect 1052 -6345 1081 -6339
rect 1623 -6343 1626 -6337
rect 1652 -6343 1655 -6317
rect 2236 -6322 2265 -6316
rect 2236 -6339 2242 -6322
rect 2259 -6323 2265 -6322
rect 2800 -6323 2803 -6317
rect 2259 -6337 2803 -6323
rect 2259 -6339 2265 -6337
rect 2236 -6345 2265 -6339
rect 2800 -6343 2803 -6337
rect 2829 -6343 2832 -6317
rect 3407 -6322 3436 -6316
rect 3407 -6339 3413 -6322
rect 3430 -6323 3436 -6322
rect 3982 -6323 3985 -6317
rect 3430 -6337 3985 -6323
rect 3430 -6339 3436 -6337
rect 3407 -6345 3436 -6339
rect 3982 -6343 3985 -6337
rect 4011 -6343 4014 -6317
rect 4594 -6322 4623 -6316
rect 4594 -6339 4600 -6322
rect 4617 -6323 4623 -6322
rect 5168 -6323 5171 -6317
rect 4617 -6337 5171 -6323
rect 4617 -6339 4623 -6337
rect 4594 -6345 4623 -6339
rect 5168 -6343 5171 -6337
rect 5197 -6343 5200 -6317
rect 5782 -6322 5811 -6316
rect 5782 -6339 5788 -6322
rect 5805 -6323 5811 -6322
rect 6347 -6323 6350 -6317
rect 5805 -6337 6350 -6323
rect 5805 -6339 5811 -6337
rect 5782 -6345 5811 -6339
rect 6347 -6343 6350 -6337
rect 6376 -6343 6379 -6317
rect 6949 -6322 6978 -6316
rect 6949 -6339 6955 -6322
rect 6972 -6323 6978 -6322
rect 7535 -6323 7538 -6317
rect 6972 -6337 7538 -6323
rect 6972 -6339 6978 -6337
rect 6949 -6345 6978 -6339
rect 7535 -6343 7538 -6337
rect 7564 -6343 7567 -6317
rect 8131 -6322 8160 -6316
rect 8131 -6339 8137 -6322
rect 8154 -6323 8160 -6322
rect 8708 -6323 8711 -6317
rect 8154 -6337 8711 -6323
rect 8154 -6339 8160 -6337
rect 8131 -6345 8160 -6339
rect 8708 -6343 8711 -6337
rect 8737 -6343 8740 -6317
rect 9317 -6322 9346 -6316
rect 9317 -6339 9323 -6322
rect 9340 -6323 9346 -6322
rect 9890 -6323 9893 -6317
rect 9340 -6337 9893 -6323
rect 9340 -6339 9346 -6337
rect 9317 -6345 9346 -6339
rect 9890 -6343 9893 -6337
rect 9919 -6343 9922 -6317
rect 10493 -6322 10522 -6316
rect 10493 -6339 10499 -6322
rect 10516 -6323 10522 -6322
rect 11079 -6323 11082 -6317
rect 10516 -6337 11082 -6323
rect 10516 -6339 10522 -6337
rect 10493 -6345 10522 -6339
rect 11079 -6343 11082 -6337
rect 11108 -6343 11111 -6317
rect 11672 -6322 11701 -6316
rect 11672 -6339 11678 -6322
rect 11695 -6323 11701 -6322
rect 12274 -6323 12277 -6317
rect 11695 -6337 12277 -6323
rect 11695 -6339 11701 -6337
rect 11672 -6345 11701 -6339
rect 12274 -6343 12277 -6337
rect 12303 -6343 12306 -6317
rect 12874 -6322 12903 -6316
rect 12874 -6339 12880 -6322
rect 12897 -6323 12903 -6322
rect 13450 -6323 13453 -6317
rect 12897 -6337 13453 -6323
rect 12897 -6339 12903 -6337
rect 12874 -6345 12903 -6339
rect 13450 -6343 13453 -6337
rect 13479 -6343 13482 -6317
rect 13773 -6322 13802 -6316
rect 13773 -6339 13779 -6322
rect 13796 -6323 13802 -6322
rect 14354 -6323 14357 -6317
rect 13796 -6337 14357 -6323
rect 13796 -6339 13802 -6337
rect 13773 -6345 13802 -6339
rect 14354 -6343 14357 -6337
rect 14383 -6343 14386 -6317
rect -4057 -6387 -4054 -6361
rect -4028 -6367 -4025 -6361
rect -4028 -6381 -3830 -6367
rect -3182 -6381 -2694 -6367
rect -2032 -6381 -1511 -6367
rect -850 -6381 -329 -6367
rect 331 -6381 852 -6367
rect 1512 -6381 2032 -6367
rect 2694 -6381 3214 -6367
rect 3876 -6381 4396 -6367
rect 5085 -6381 5578 -6367
rect 6240 -6381 6760 -6367
rect 7422 -6381 7942 -6367
rect 8604 -6381 9126 -6367
rect 9788 -6381 10310 -6367
rect 10972 -6381 11497 -6367
rect 12159 -6381 12684 -6367
rect 13346 -6381 13585 -6367
rect -4028 -6387 -4025 -6381
rect -4123 -6427 -4120 -6401
rect -4094 -6407 -4091 -6401
rect -4094 -6421 -3829 -6407
rect -3182 -6421 -2694 -6407
rect -2032 -6421 -1511 -6407
rect -850 -6421 -329 -6407
rect 331 -6421 852 -6407
rect 1512 -6421 2032 -6407
rect 2694 -6421 3214 -6407
rect 3876 -6421 4396 -6407
rect 5085 -6421 5578 -6407
rect 6240 -6421 6760 -6407
rect 7422 -6421 7942 -6407
rect 8604 -6421 9126 -6407
rect 9788 -6421 10310 -6407
rect 10972 -6421 11497 -6407
rect 12159 -6421 12684 -6407
rect 13346 -6421 13585 -6407
rect -4094 -6427 -4091 -6421
rect -3916 -7105 -3913 -7079
rect -3887 -7085 -3884 -7079
rect -3887 -7099 -3830 -7085
rect -3196 -7099 -2694 -7085
rect -2046 -7099 -1512 -7085
rect -864 -7099 -330 -7085
rect 317 -7099 850 -7085
rect 1498 -7099 2032 -7085
rect 2680 -7099 3214 -7085
rect 3862 -7099 4396 -7085
rect 5044 -7099 5578 -7085
rect 6226 -7099 6760 -7085
rect 7408 -7099 7943 -7085
rect 8590 -7099 9126 -7085
rect 9774 -7099 10311 -7085
rect 10957 -7099 11501 -7085
rect 12145 -7099 12684 -7085
rect 13332 -7099 13585 -7085
rect -3887 -7105 -3884 -7099
rect -3221 -7176 -3192 -7174
rect -2071 -7176 -2042 -7173
rect -889 -7176 -860 -7173
rect 292 -7176 321 -7173
rect 1473 -7176 1502 -7173
rect 2655 -7176 2684 -7173
rect 3837 -7176 3866 -7173
rect 5019 -7176 5048 -7173
rect 6201 -7176 6230 -7173
rect 7383 -7176 7412 -7173
rect 8565 -7176 8594 -7173
rect 9749 -7176 9778 -7173
rect 10933 -7176 10962 -7173
rect 12120 -7176 12149 -7173
rect 13307 -7176 13336 -7173
rect 14208 -7176 14237 -7173
rect 14553 -7176 14556 -7171
rect -3221 -7177 -2065 -7176
rect -3221 -7194 -3215 -7177
rect -3198 -7193 -2065 -7177
rect -2048 -7193 -883 -7176
rect -866 -7193 298 -7176
rect 315 -7193 1479 -7176
rect 1496 -7193 2661 -7176
rect 2678 -7193 3843 -7176
rect 3860 -7193 5025 -7176
rect 5042 -7193 6207 -7176
rect 6224 -7193 7389 -7176
rect 7406 -7193 8571 -7176
rect 8588 -7193 9755 -7176
rect 9772 -7193 10939 -7176
rect 10956 -7193 12126 -7176
rect 12143 -7193 13313 -7176
rect 13330 -7193 14214 -7176
rect 14231 -7193 14556 -7176
rect -3198 -7194 -3192 -7193
rect -3221 -7197 -3192 -7194
rect -2071 -7196 -2042 -7193
rect -889 -7196 -860 -7193
rect 292 -7196 321 -7193
rect 1473 -7196 1502 -7193
rect 2655 -7196 2684 -7193
rect 3837 -7196 3866 -7193
rect 5019 -7196 5048 -7193
rect 6201 -7196 6230 -7193
rect 7383 -7196 7412 -7193
rect 8565 -7196 8594 -7193
rect 9749 -7196 9778 -7193
rect 10933 -7196 10962 -7193
rect 12120 -7196 12149 -7193
rect 13307 -7196 13336 -7193
rect 14208 -7196 14237 -7193
rect 14553 -7197 14556 -7193
rect 14582 -7197 14585 -7171
rect -3221 -7273 -3192 -7271
rect -2071 -7273 -2042 -7270
rect -889 -7273 -860 -7270
rect 292 -7273 321 -7270
rect 1473 -7273 1502 -7270
rect 2655 -7273 2684 -7270
rect 3837 -7273 3866 -7270
rect 5019 -7273 5048 -7270
rect 6201 -7273 6230 -7270
rect 7383 -7273 7412 -7270
rect 8565 -7273 8594 -7270
rect 9749 -7273 9778 -7270
rect 10933 -7273 10962 -7270
rect 12120 -7273 12149 -7270
rect 13307 -7273 13336 -7270
rect 14211 -7273 14234 -7267
rect 14608 -7273 14611 -7268
rect -3221 -7274 -2065 -7273
rect -3221 -7291 -3215 -7274
rect -3198 -7290 -2065 -7274
rect -2048 -7290 -883 -7273
rect -866 -7290 298 -7273
rect 315 -7290 1479 -7273
rect 1496 -7290 2661 -7273
rect 2678 -7290 3843 -7273
rect 3860 -7290 5025 -7273
rect 5042 -7290 6207 -7273
rect 6224 -7290 7389 -7273
rect 7406 -7290 8571 -7273
rect 8588 -7290 9755 -7273
rect 9772 -7290 10939 -7273
rect 10956 -7290 12126 -7273
rect 12143 -7290 13313 -7273
rect 13330 -7290 14214 -7273
rect 14231 -7290 14611 -7273
rect -3198 -7291 -3192 -7290
rect -3221 -7294 -3192 -7291
rect -2071 -7293 -2042 -7290
rect -889 -7293 -860 -7290
rect 292 -7293 321 -7290
rect 1473 -7293 1502 -7290
rect 2655 -7293 2684 -7290
rect 3837 -7293 3866 -7290
rect 5019 -7293 5048 -7290
rect 6201 -7293 6230 -7290
rect 7383 -7293 7412 -7290
rect 8565 -7293 8594 -7290
rect 9749 -7293 9778 -7290
rect 10933 -7293 10962 -7290
rect 12120 -7293 12149 -7290
rect 13307 -7293 13336 -7290
rect 14211 -7296 14234 -7290
rect 14608 -7294 14611 -7290
rect 14637 -7294 14640 -7268
rect -3913 -7369 -3887 -7366
rect -3887 -7389 -3844 -7375
rect -3196 -7389 -2694 -7375
rect -2046 -7389 -1512 -7375
rect -864 -7389 -331 -7375
rect 317 -7389 850 -7375
rect 1498 -7389 2033 -7375
rect 2680 -7389 3216 -7375
rect 3862 -7389 4397 -7375
rect 5044 -7389 5578 -7375
rect 6226 -7389 6760 -7375
rect 7408 -7389 7942 -7375
rect 8590 -7389 9126 -7375
rect 9774 -7389 10310 -7375
rect 10958 -7389 11497 -7375
rect 12145 -7389 12684 -7375
rect 13332 -7389 13585 -7375
rect -3913 -7398 -3887 -7395
rect -4123 -8073 -4120 -8047
rect -4094 -8053 -4091 -8047
rect -4094 -8067 -3826 -8053
rect -3196 -8067 -2694 -8053
rect -2046 -8067 -1512 -8053
rect -864 -8067 -330 -8053
rect 317 -8067 850 -8053
rect 1498 -8067 2033 -8053
rect 2680 -8067 3215 -8053
rect 3862 -8067 4396 -8053
rect 5044 -8067 5578 -8053
rect 6224 -8067 6760 -8053
rect 7408 -8067 7943 -8053
rect 8590 -8067 9127 -8053
rect 9774 -8067 10311 -8053
rect 10956 -8067 11498 -8053
rect 12145 -8067 12684 -8053
rect 13332 -8067 13586 -8053
rect -4094 -8073 -4091 -8067
rect -4057 -8113 -4054 -8087
rect -4028 -8093 -4025 -8087
rect -4028 -8107 -3830 -8093
rect -3182 -8107 -2680 -8093
rect -2032 -8107 -1497 -8093
rect -850 -8107 -317 -8093
rect 331 -8107 864 -8093
rect 1502 -8107 2046 -8093
rect 2689 -8107 3228 -8093
rect 3875 -8107 4410 -8093
rect 5057 -8107 5592 -8093
rect 6240 -8107 6774 -8093
rect 7421 -8107 7956 -8093
rect 8604 -8107 9140 -8093
rect 9784 -8107 10324 -8093
rect 10967 -8107 11511 -8093
rect 12159 -8107 12698 -8093
rect 13346 -8107 13599 -8093
rect -4028 -8113 -4025 -8107
rect -3646 -8135 -3623 -8129
rect -3646 -8152 -3643 -8135
rect -3626 -8136 -3623 -8135
rect -3029 -8136 -3026 -8130
rect -3626 -8150 -3026 -8136
rect -3626 -8152 -3623 -8150
rect -3646 -8158 -3623 -8152
rect -3029 -8156 -3026 -8150
rect -3000 -8156 -2997 -8130
rect -2514 -8135 -2485 -8129
rect -2514 -8152 -2508 -8135
rect -2491 -8136 -2485 -8135
rect -1873 -8136 -1870 -8130
rect -2491 -8150 -1870 -8136
rect -2491 -8152 -2485 -8150
rect -2514 -8158 -2485 -8152
rect -1873 -8156 -1870 -8150
rect -1844 -8156 -1841 -8130
rect -1339 -8135 -1310 -8129
rect -1339 -8152 -1333 -8135
rect -1316 -8136 -1310 -8135
rect -704 -8136 -701 -8130
rect -1316 -8150 -701 -8136
rect -1316 -8152 -1310 -8150
rect -1339 -8158 -1310 -8152
rect -704 -8156 -701 -8150
rect -675 -8156 -672 -8130
rect -157 -8135 -128 -8129
rect -157 -8152 -151 -8135
rect -134 -8136 -128 -8135
rect 487 -8136 490 -8130
rect -134 -8150 490 -8136
rect -134 -8152 -128 -8150
rect -157 -8158 -128 -8152
rect 487 -8156 490 -8150
rect 516 -8156 519 -8130
rect 1025 -8135 1054 -8129
rect 1025 -8152 1031 -8135
rect 1048 -8136 1054 -8135
rect 1664 -8136 1667 -8130
rect 1048 -8150 1667 -8136
rect 1048 -8152 1054 -8150
rect 1025 -8158 1054 -8152
rect 1664 -8156 1667 -8150
rect 1693 -8156 1696 -8130
rect 2207 -8135 2236 -8129
rect 2207 -8152 2213 -8135
rect 2230 -8136 2236 -8135
rect 2841 -8136 2844 -8130
rect 2230 -8150 2844 -8136
rect 2230 -8152 2236 -8150
rect 2207 -8158 2236 -8152
rect 2841 -8156 2844 -8150
rect 2870 -8156 2873 -8130
rect 3401 -8135 3430 -8129
rect 3401 -8152 3407 -8135
rect 3424 -8136 3430 -8135
rect 4023 -8136 4026 -8130
rect 3424 -8150 4026 -8136
rect 3424 -8152 3430 -8150
rect 3401 -8158 3430 -8152
rect 4023 -8156 4026 -8150
rect 4052 -8156 4055 -8130
rect 4578 -8135 4607 -8129
rect 4578 -8152 4584 -8135
rect 4601 -8136 4607 -8135
rect 5209 -8136 5212 -8130
rect 4601 -8150 5212 -8136
rect 4601 -8152 4607 -8150
rect 4578 -8158 4607 -8152
rect 5209 -8156 5212 -8150
rect 5238 -8156 5241 -8130
rect 5761 -8135 5790 -8129
rect 5761 -8152 5767 -8135
rect 5784 -8136 5790 -8135
rect 6388 -8136 6391 -8130
rect 5784 -8150 6391 -8136
rect 5784 -8152 5790 -8150
rect 5761 -8158 5790 -8152
rect 6388 -8156 6391 -8150
rect 6417 -8156 6420 -8130
rect 6934 -8135 6963 -8129
rect 6934 -8152 6940 -8135
rect 6957 -8136 6963 -8135
rect 7576 -8136 7579 -8130
rect 6957 -8150 7579 -8136
rect 6957 -8152 6963 -8150
rect 6934 -8158 6963 -8152
rect 7576 -8156 7579 -8150
rect 7605 -8156 7608 -8130
rect 8117 -8135 8146 -8129
rect 8117 -8152 8123 -8135
rect 8140 -8136 8146 -8135
rect 8749 -8136 8752 -8130
rect 8140 -8150 8752 -8136
rect 8140 -8152 8146 -8150
rect 8117 -8158 8146 -8152
rect 8749 -8156 8752 -8150
rect 8778 -8156 8781 -8130
rect 9300 -8135 9329 -8129
rect 9300 -8152 9306 -8135
rect 9323 -8136 9329 -8135
rect 9931 -8136 9934 -8130
rect 9323 -8150 9934 -8136
rect 9323 -8152 9329 -8150
rect 9300 -8158 9329 -8152
rect 9931 -8156 9934 -8150
rect 9960 -8156 9963 -8130
rect 10478 -8135 10507 -8129
rect 10478 -8152 10484 -8135
rect 10501 -8136 10507 -8135
rect 11120 -8136 11123 -8130
rect 10501 -8150 11123 -8136
rect 10501 -8152 10507 -8150
rect 10478 -8158 10507 -8152
rect 11120 -8156 11123 -8150
rect 11149 -8156 11152 -8130
rect 11672 -8135 11701 -8129
rect 11672 -8152 11678 -8135
rect 11695 -8136 11701 -8135
rect 12315 -8136 12318 -8130
rect 11695 -8150 12318 -8136
rect 11695 -8152 11701 -8150
rect 11672 -8158 11701 -8152
rect 12315 -8156 12318 -8150
rect 12344 -8156 12347 -8130
rect 12867 -8135 12896 -8129
rect 12867 -8152 12873 -8135
rect 12890 -8136 12896 -8135
rect 13491 -8136 13494 -8130
rect 12890 -8150 13494 -8136
rect 12890 -8152 12896 -8150
rect 12867 -8158 12896 -8152
rect 13491 -8156 13494 -8150
rect 13520 -8156 13523 -8130
rect 13772 -8135 13801 -8129
rect 13772 -8152 13778 -8135
rect 13795 -8136 13801 -8135
rect 14395 -8136 14398 -8130
rect 13795 -8150 14398 -8136
rect 13795 -8152 13801 -8150
rect 13772 -8158 13801 -8152
rect 14395 -8156 14398 -8150
rect 14424 -8156 14427 -8130
rect -3991 -8616 -3988 -8590
rect -3962 -8596 -3959 -8590
rect -3962 -8610 -3844 -8596
rect -3196 -8610 -2694 -8596
rect -2046 -8610 -1512 -8596
rect -864 -8610 -330 -8596
rect 317 -8610 850 -8596
rect 1498 -8610 2032 -8596
rect 2680 -8610 3214 -8596
rect 3862 -8610 4396 -8596
rect 5044 -8610 5578 -8596
rect 6226 -8610 6760 -8596
rect 7407 -8610 7942 -8596
rect 8590 -8610 9128 -8596
rect 9772 -8610 10310 -8596
rect 10958 -8610 11497 -8596
rect 12145 -8610 12684 -8596
rect 13332 -8610 13585 -8596
rect -3962 -8616 -3959 -8610
<< via1 >>
rect 129 4838 155 4864
rect 128 4755 154 4781
rect 130 4669 156 4695
rect 128 4597 154 4623
rect 129 4512 155 4538
rect 129 4432 155 4458
rect 128 4356 154 4382
rect 130 4219 156 4245
rect 130 4133 156 4159
rect 128 4059 154 4085
rect 130 3976 156 4002
rect 130 3892 156 3918
rect 129 3818 155 3844
rect 129 3577 155 3603
rect 129 3336 155 3362
rect 129 3095 155 3121
rect 129 2854 155 2880
rect 128 2573 154 2599
rect 129 2332 155 2358
rect 129 2091 155 2117
rect 129 1850 155 1876
rect 129 1609 155 1635
rect 129 1368 155 1394
rect 128 1127 154 1153
rect 129 886 155 912
rect 128 604 154 630
rect 130 363 156 389
rect 129 122 155 148
rect 129 -119 155 -93
rect 129 -204 155 -178
rect 129 -283 155 -257
rect 129 -360 155 -334
rect 129 -442 155 -416
rect 130 -521 156 -495
rect 129 -601 155 -575
rect 129 -744 155 -718
rect 129 -824 155 -798
rect 129 -901 155 -875
rect 129 -981 155 -955
rect 130 -1068 156 -1042
rect 129 -1142 155 -1116
rect 597 -1391 623 -1386
rect 597 -1408 601 -1391
rect 601 -1408 618 -1391
rect 618 -1408 623 -1391
rect 597 -1412 623 -1408
rect 1172 -1392 1198 -1387
rect 1172 -1409 1176 -1392
rect 1176 -1409 1193 -1392
rect 1193 -1409 1198 -1392
rect 1172 -1413 1198 -1409
rect 1747 -1394 1773 -1389
rect 1747 -1411 1751 -1394
rect 1751 -1411 1768 -1394
rect 1768 -1411 1773 -1394
rect 1747 -1415 1773 -1411
rect 2322 -1394 2348 -1389
rect 2322 -1411 2326 -1394
rect 2326 -1411 2343 -1394
rect 2343 -1411 2348 -1394
rect 2322 -1415 2348 -1411
rect 2897 -1392 2923 -1387
rect 2897 -1409 2901 -1392
rect 2901 -1409 2918 -1392
rect 2918 -1409 2923 -1392
rect 2897 -1413 2923 -1409
rect 3472 -1389 3498 -1384
rect 3472 -1406 3476 -1389
rect 3476 -1406 3493 -1389
rect 3493 -1406 3498 -1389
rect 3472 -1410 3498 -1406
rect 4047 -1387 4073 -1382
rect 4047 -1404 4051 -1387
rect 4051 -1404 4068 -1387
rect 4068 -1404 4073 -1387
rect 4047 -1408 4073 -1404
rect 4622 -1387 4648 -1382
rect 4622 -1404 4626 -1387
rect 4626 -1404 4643 -1387
rect 4643 -1404 4648 -1387
rect 4622 -1408 4648 -1404
rect 5197 -1392 5223 -1387
rect 5197 -1409 5201 -1392
rect 5201 -1409 5218 -1392
rect 5218 -1409 5223 -1392
rect 5197 -1413 5223 -1409
rect 5772 -1389 5798 -1384
rect 5772 -1406 5776 -1389
rect 5776 -1406 5793 -1389
rect 5793 -1406 5798 -1389
rect 5772 -1410 5798 -1406
rect 6347 -1393 6373 -1388
rect 6347 -1410 6351 -1393
rect 6351 -1410 6368 -1393
rect 6368 -1410 6373 -1393
rect 6347 -1414 6373 -1410
rect 6922 -1394 6948 -1389
rect 6922 -1411 6926 -1394
rect 6926 -1411 6943 -1394
rect 6943 -1411 6948 -1394
rect 6922 -1415 6948 -1411
rect 7497 -1390 7523 -1385
rect 7497 -1407 7501 -1390
rect 7501 -1407 7518 -1390
rect 7518 -1407 7523 -1390
rect 7497 -1411 7523 -1407
rect 8072 -1394 8098 -1389
rect 8072 -1411 8076 -1394
rect 8076 -1411 8093 -1394
rect 8093 -1411 8098 -1394
rect 8072 -1415 8098 -1411
rect 8647 -1390 8673 -1385
rect 8647 -1407 8651 -1390
rect 8651 -1407 8668 -1390
rect 8668 -1407 8673 -1390
rect 8647 -1411 8673 -1407
rect 9222 -1391 9248 -1386
rect 9222 -1408 9226 -1391
rect 9226 -1408 9243 -1391
rect 9243 -1408 9248 -1391
rect 9222 -1412 9248 -1408
rect 129 -1919 155 -1893
rect -33 -2058 -7 -2032
rect 130 -2059 156 -2033
rect 228 -2127 254 -2101
rect 809 -2125 835 -2099
rect 1381 -2126 1407 -2100
rect 1959 -2128 1985 -2102
rect 2534 -2128 2560 -2102
rect 3105 -2130 3131 -2104
rect 3682 -2129 3708 -2103
rect 4262 -2128 4288 -2102
rect 4832 -2127 4858 -2101
rect 5409 -2129 5435 -2103
rect 5983 -2127 6009 -2101
rect 6556 -2128 6582 -2102
rect 7133 -2129 7159 -2103
rect 7709 -2129 7735 -2103
rect 8282 -2131 8308 -2105
rect 8857 -2131 8883 -2105
rect 299 -2300 325 -2274
rect 752 -2300 778 -2274
rect 874 -2300 900 -2274
rect 1327 -2300 1353 -2274
rect 1449 -2300 1475 -2274
rect 1902 -2300 1928 -2274
rect 2024 -2300 2050 -2274
rect 2477 -2300 2503 -2274
rect 2599 -2300 2625 -2274
rect 3052 -2300 3078 -2274
rect 3174 -2300 3200 -2274
rect 3627 -2300 3653 -2274
rect 3749 -2300 3775 -2274
rect 4202 -2300 4228 -2274
rect 4324 -2300 4350 -2274
rect 4777 -2300 4803 -2274
rect 4899 -2300 4925 -2274
rect 5352 -2300 5378 -2274
rect 5474 -2300 5500 -2274
rect 5927 -2300 5953 -2274
rect 6049 -2300 6075 -2274
rect 6502 -2300 6528 -2274
rect 6624 -2300 6650 -2274
rect 7077 -2300 7103 -2274
rect 7199 -2300 7225 -2274
rect 7652 -2300 7678 -2274
rect 7774 -2300 7800 -2274
rect 8227 -2300 8253 -2274
rect 8349 -2300 8375 -2274
rect 8802 -2300 8828 -2274
rect 8924 -2300 8950 -2274
rect 9377 -2300 9403 -2274
rect 526 -2344 552 -2341
rect 526 -2364 529 -2344
rect 529 -2364 549 -2344
rect 549 -2364 552 -2344
rect 526 -2367 552 -2364
rect 813 -2327 839 -2322
rect 813 -2344 817 -2327
rect 817 -2344 834 -2327
rect 834 -2344 839 -2327
rect 813 -2348 839 -2344
rect 1101 -2345 1127 -2342
rect 1101 -2365 1104 -2345
rect 1104 -2365 1124 -2345
rect 1124 -2365 1127 -2345
rect 1101 -2368 1127 -2365
rect 1676 -2350 1702 -2347
rect 1676 -2370 1679 -2350
rect 1679 -2370 1699 -2350
rect 1699 -2370 1702 -2350
rect 1676 -2373 1702 -2370
rect 1962 -2328 1988 -2323
rect 1962 -2345 1966 -2328
rect 1966 -2345 1983 -2328
rect 1983 -2345 1988 -2328
rect 1962 -2349 1988 -2345
rect 2251 -2350 2277 -2347
rect 2251 -2370 2254 -2350
rect 2254 -2370 2274 -2350
rect 2274 -2370 2277 -2350
rect 2251 -2373 2277 -2370
rect 2826 -2350 2852 -2347
rect 2826 -2370 2829 -2350
rect 2829 -2370 2849 -2350
rect 2849 -2370 2852 -2350
rect 2826 -2373 2852 -2370
rect 3105 -2329 3131 -2324
rect 3105 -2346 3109 -2329
rect 3109 -2346 3126 -2329
rect 3126 -2346 3131 -2329
rect 3105 -2350 3131 -2346
rect 3401 -2350 3427 -2347
rect 3401 -2370 3404 -2350
rect 3404 -2370 3424 -2350
rect 3424 -2370 3427 -2350
rect 3401 -2373 3427 -2370
rect 3976 -2350 4002 -2347
rect 3976 -2370 3979 -2350
rect 3979 -2370 3999 -2350
rect 3999 -2370 4002 -2350
rect 3976 -2373 4002 -2370
rect 4262 -2330 4288 -2325
rect 4262 -2347 4266 -2330
rect 4266 -2347 4283 -2330
rect 4283 -2347 4288 -2330
rect 4262 -2351 4288 -2347
rect 4551 -2350 4577 -2347
rect 4551 -2370 4554 -2350
rect 4554 -2370 4574 -2350
rect 4574 -2370 4577 -2350
rect 4551 -2373 4577 -2370
rect 5126 -2350 5152 -2347
rect 5126 -2370 5129 -2350
rect 5129 -2370 5149 -2350
rect 5149 -2370 5152 -2350
rect 5126 -2373 5152 -2370
rect 5402 -2328 5428 -2323
rect 5402 -2345 5406 -2328
rect 5406 -2345 5423 -2328
rect 5423 -2345 5428 -2328
rect 5402 -2349 5428 -2345
rect 5701 -2350 5727 -2347
rect 5701 -2370 5704 -2350
rect 5704 -2370 5724 -2350
rect 5724 -2370 5727 -2350
rect 5701 -2373 5727 -2370
rect 6276 -2350 6302 -2347
rect 6276 -2370 6279 -2350
rect 6279 -2370 6299 -2350
rect 6299 -2370 6302 -2350
rect 6276 -2373 6302 -2370
rect 6570 -2328 6596 -2323
rect 6570 -2345 6574 -2328
rect 6574 -2345 6591 -2328
rect 6591 -2345 6596 -2328
rect 6570 -2349 6596 -2345
rect 6851 -2350 6877 -2347
rect 6851 -2370 6854 -2350
rect 6854 -2370 6874 -2350
rect 6874 -2370 6877 -2350
rect 6851 -2373 6877 -2370
rect 7426 -2350 7452 -2347
rect 7426 -2370 7429 -2350
rect 7429 -2370 7449 -2350
rect 7449 -2370 7452 -2350
rect 7426 -2373 7452 -2370
rect 7715 -2328 7741 -2323
rect 7715 -2345 7719 -2328
rect 7719 -2345 7736 -2328
rect 7736 -2345 7741 -2328
rect 7715 -2349 7741 -2345
rect 8872 -2326 8898 -2321
rect 8872 -2343 8876 -2326
rect 8876 -2343 8893 -2326
rect 8893 -2343 8898 -2326
rect 8872 -2347 8898 -2343
rect 8001 -2350 8027 -2347
rect 8001 -2370 8004 -2350
rect 8004 -2370 8024 -2350
rect 8024 -2370 8027 -2350
rect 8001 -2373 8027 -2370
rect 8576 -2350 8602 -2347
rect 8576 -2370 8579 -2350
rect 8579 -2370 8599 -2350
rect 8599 -2370 8602 -2350
rect 8576 -2373 8602 -2370
rect 9151 -2350 9177 -2347
rect 9151 -2370 9154 -2350
rect 9154 -2370 9174 -2350
rect 9174 -2370 9177 -2350
rect 9151 -2373 9177 -2370
rect 737 -2426 763 -2421
rect 737 -2443 741 -2426
rect 741 -2443 758 -2426
rect 758 -2443 763 -2426
rect 737 -2447 763 -2443
rect 892 -2426 918 -2421
rect 892 -2443 896 -2426
rect 896 -2443 913 -2426
rect 913 -2443 918 -2426
rect 892 -2447 918 -2443
rect 1887 -2426 1913 -2421
rect 1887 -2443 1891 -2426
rect 1891 -2443 1908 -2426
rect 1908 -2443 1913 -2426
rect 1887 -2447 1913 -2443
rect 2042 -2426 2068 -2421
rect 2042 -2443 2046 -2426
rect 2046 -2443 2063 -2426
rect 2063 -2443 2068 -2426
rect 2042 -2447 2068 -2443
rect 3037 -2426 3063 -2421
rect 3037 -2443 3041 -2426
rect 3041 -2443 3058 -2426
rect 3058 -2443 3063 -2426
rect 3037 -2447 3063 -2443
rect 3191 -2426 3217 -2421
rect 3191 -2443 3195 -2426
rect 3195 -2443 3212 -2426
rect 3212 -2443 3217 -2426
rect 3191 -2447 3217 -2443
rect 4184 -2426 4210 -2421
rect 4184 -2443 4188 -2426
rect 4188 -2443 4205 -2426
rect 4205 -2443 4210 -2426
rect 4184 -2447 4210 -2443
rect 4343 -2427 4369 -2422
rect 4343 -2444 4347 -2427
rect 4347 -2444 4364 -2427
rect 4364 -2444 4369 -2427
rect 4343 -2448 4369 -2444
rect -3924 -2484 -3898 -2458
rect 5336 -2426 5362 -2421
rect 5336 -2443 5340 -2426
rect 5340 -2443 5357 -2426
rect 5357 -2443 5362 -2426
rect 5336 -2447 5362 -2443
rect 5491 -2426 5517 -2421
rect 5491 -2443 5495 -2426
rect 5495 -2443 5512 -2426
rect 5512 -2443 5517 -2426
rect 5491 -2447 5517 -2443
rect 6487 -2427 6513 -2422
rect 6487 -2444 6491 -2427
rect 6491 -2444 6508 -2427
rect 6508 -2444 6513 -2427
rect 6487 -2448 6513 -2444
rect 6640 -2427 6666 -2422
rect 6640 -2444 6644 -2427
rect 6644 -2444 6661 -2427
rect 6661 -2444 6666 -2427
rect 6640 -2448 6666 -2444
rect 7638 -2426 7664 -2421
rect 7638 -2443 7642 -2426
rect 7642 -2443 7659 -2426
rect 7659 -2443 7664 -2426
rect 7638 -2447 7664 -2443
rect 7791 -2426 7817 -2421
rect 7791 -2443 7795 -2426
rect 7795 -2443 7812 -2426
rect 7812 -2443 7817 -2426
rect 7791 -2447 7817 -2443
rect 8787 -2425 8813 -2420
rect 8787 -2442 8791 -2425
rect 8791 -2442 8808 -2425
rect 8808 -2442 8813 -2425
rect 8787 -2446 8813 -2442
rect 8939 -2426 8965 -2421
rect 8939 -2443 8943 -2426
rect 8943 -2443 8960 -2426
rect 8960 -2443 8965 -2426
rect 8939 -2447 8965 -2443
rect 468 -2503 494 -2498
rect 468 -2520 472 -2503
rect 472 -2520 489 -2503
rect 489 -2520 494 -2503
rect 468 -2524 494 -2520
rect 1161 -2496 1187 -2491
rect 1161 -2513 1165 -2496
rect 1165 -2513 1182 -2496
rect 1182 -2513 1187 -2496
rect 1161 -2517 1187 -2513
rect 1617 -2495 1643 -2490
rect 1617 -2512 1621 -2495
rect 1621 -2512 1638 -2495
rect 1638 -2512 1643 -2495
rect 1617 -2516 1643 -2512
rect 2310 -2500 2336 -2495
rect 2310 -2517 2314 -2500
rect 2314 -2517 2331 -2500
rect 2331 -2517 2336 -2500
rect 2310 -2521 2336 -2517
rect 2769 -2501 2795 -2496
rect 2769 -2518 2773 -2501
rect 2773 -2518 2790 -2501
rect 2790 -2518 2795 -2501
rect 2769 -2522 2795 -2518
rect 3461 -2499 3487 -2494
rect 3461 -2516 3465 -2499
rect 3465 -2516 3482 -2499
rect 3482 -2516 3487 -2499
rect 3461 -2520 3487 -2516
rect 3919 -2501 3945 -2496
rect 3919 -2518 3923 -2501
rect 3923 -2518 3940 -2501
rect 3940 -2518 3945 -2501
rect 3919 -2522 3945 -2518
rect 4610 -2503 4636 -2498
rect 4610 -2520 4614 -2503
rect 4614 -2520 4631 -2503
rect 4631 -2520 4636 -2503
rect 4610 -2524 4636 -2520
rect 5068 -2497 5094 -2492
rect 5068 -2514 5072 -2497
rect 5072 -2514 5089 -2497
rect 5089 -2514 5094 -2497
rect 5068 -2518 5094 -2514
rect 5761 -2499 5787 -2494
rect 5761 -2516 5765 -2499
rect 5765 -2516 5782 -2499
rect 5782 -2516 5787 -2499
rect 5761 -2520 5787 -2516
rect 6218 -2495 6244 -2490
rect 6218 -2512 6222 -2495
rect 6222 -2512 6239 -2495
rect 6239 -2512 6244 -2495
rect 6218 -2516 6244 -2512
rect 6910 -2499 6936 -2494
rect 6910 -2516 6914 -2499
rect 6914 -2516 6931 -2499
rect 6931 -2516 6936 -2499
rect 6910 -2520 6936 -2516
rect 7368 -2499 7394 -2494
rect 7368 -2516 7372 -2499
rect 7372 -2516 7389 -2499
rect 7389 -2516 7394 -2499
rect 7368 -2520 7394 -2516
rect 8060 -2502 8086 -2497
rect 8060 -2519 8064 -2502
rect 8064 -2519 8081 -2502
rect 8081 -2519 8086 -2502
rect 8060 -2523 8086 -2519
rect 8518 -2500 8544 -2495
rect 8518 -2517 8522 -2500
rect 8522 -2517 8539 -2500
rect 8539 -2517 8544 -2500
rect 8518 -2521 8544 -2517
rect 9206 -2494 9236 -2491
rect 9206 -2518 9209 -2494
rect 9209 -2518 9233 -2494
rect 9233 -2518 9236 -2494
rect 9206 -2521 9236 -2518
rect -2744 -2566 -2718 -2540
rect 13532 -2563 13558 -2537
rect -1565 -2629 -1539 -2603
rect 12586 -2613 12612 -2587
rect 11423 -2663 11449 -2637
rect -387 -2704 -361 -2678
rect 10210 -2726 10236 -2700
rect 811 -2775 837 -2749
rect 9036 -2789 9062 -2763
rect 1978 -2855 2004 -2829
rect 7848 -2861 7874 -2835
rect 3137 -2939 3163 -2913
rect 6646 -2941 6672 -2915
rect 4311 -3010 4337 -2984
rect 5496 -3028 5522 -3002
rect -3988 -3151 -3962 -3125
rect -3148 -3610 -3122 -3584
rect -1993 -3610 -1967 -3584
rect -824 -3610 -798 -3584
rect 367 -3610 393 -3584
rect 1544 -3610 1570 -3584
rect 2721 -3610 2747 -3584
rect 3903 -3610 3929 -3584
rect 5089 -3610 5115 -3584
rect 6268 -3610 6294 -3584
rect 7456 -3610 7482 -3584
rect 8629 -3610 8655 -3584
rect 9811 -3610 9837 -3584
rect 11000 -3610 11026 -3584
rect 12195 -3610 12221 -3584
rect 13371 -3610 13397 -3584
rect 14275 -3610 14301 -3584
rect -4054 -3654 -4028 -3628
rect -4120 -3694 -4094 -3668
rect -3927 -4163 -3895 -4131
rect -2743 -4161 -2717 -4135
rect -1564 -4161 -1538 -4135
rect -386 -4161 -360 -4135
rect 812 -4161 838 -4135
rect 1979 -4160 2005 -4134
rect 3138 -4159 3164 -4133
rect 4312 -4159 4338 -4133
rect 5497 -4159 5523 -4133
rect 6647 -4161 6673 -4135
rect 7849 -4161 7875 -4135
rect 9037 -4161 9063 -4135
rect 10211 -4161 10237 -4135
rect 11424 -4160 11450 -4134
rect 12587 -4161 12613 -4135
rect 13533 -4160 13559 -4134
rect -4178 -4372 -4152 -4346
rect -3913 -4372 -3887 -4346
rect 14446 -4471 14472 -4445
rect 14502 -4560 14528 -4534
rect -3913 -4662 -3887 -4636
rect -4120 -5340 -4094 -5314
rect -4054 -5380 -4028 -5354
rect -3107 -5423 -3081 -5397
rect -1953 -5423 -1927 -5397
rect -784 -5423 -758 -5397
rect 407 -5423 433 -5397
rect 1584 -5423 1610 -5397
rect 2761 -5423 2787 -5397
rect 3943 -5423 3969 -5397
rect 5129 -5423 5155 -5397
rect 6308 -5423 6334 -5397
rect 7496 -5423 7522 -5397
rect 8669 -5423 8695 -5397
rect 9851 -5423 9877 -5397
rect 11040 -5423 11066 -5397
rect 12235 -5423 12261 -5397
rect 13411 -5423 13437 -5397
rect 14315 -5423 14341 -5397
rect -3987 -5883 -3961 -5857
rect -3067 -6343 -3041 -6317
rect -1911 -6343 -1885 -6317
rect -742 -6343 -716 -6317
rect 449 -6343 475 -6317
rect 1626 -6343 1652 -6317
rect 2803 -6343 2829 -6317
rect 3985 -6343 4011 -6317
rect 5171 -6343 5197 -6317
rect 6350 -6343 6376 -6317
rect 7538 -6343 7564 -6317
rect 8711 -6343 8737 -6317
rect 9893 -6343 9919 -6317
rect 11082 -6343 11108 -6317
rect 12277 -6343 12303 -6317
rect 13453 -6343 13479 -6317
rect 14357 -6343 14383 -6317
rect -4054 -6387 -4028 -6361
rect -4120 -6427 -4094 -6401
rect -3913 -7105 -3887 -7079
rect 14556 -7197 14582 -7171
rect 14611 -7294 14637 -7268
rect -3913 -7395 -3887 -7369
rect -4120 -8073 -4094 -8047
rect -4054 -8113 -4028 -8087
rect -3026 -8156 -3000 -8130
rect -1870 -8156 -1844 -8130
rect -701 -8156 -675 -8130
rect 490 -8156 516 -8130
rect 1667 -8156 1693 -8130
rect 2844 -8156 2870 -8130
rect 4026 -8156 4052 -8130
rect 5212 -8156 5238 -8130
rect 6391 -8156 6417 -8130
rect 7579 -8156 7605 -8130
rect 8752 -8156 8778 -8130
rect 9934 -8156 9960 -8130
rect 11123 -8156 11149 -8130
rect 12318 -8156 12344 -8130
rect 13494 -8156 13520 -8130
rect 14398 -8156 14424 -8130
rect -3988 -8616 -3962 -8590
<< metal2 >>
rect -4314 5061 -4284 5066
rect -4314 5026 -4284 5031
rect -4306 -3058 -4292 5026
rect 129 4864 155 4867
rect 129 4835 155 4838
rect 135 4784 150 4835
rect 125 4781 157 4784
rect 125 4755 128 4781
rect 154 4755 157 4781
rect 125 4752 157 4755
rect 135 4698 150 4752
rect 127 4695 159 4698
rect 127 4669 130 4695
rect 156 4669 159 4695
rect 127 4666 159 4669
rect 135 4626 150 4666
rect 128 4623 154 4626
rect 128 4594 154 4597
rect 135 4541 150 4594
rect 126 4538 158 4541
rect 126 4512 129 4538
rect 155 4512 158 4538
rect 126 4509 158 4512
rect 135 4461 150 4509
rect 126 4458 158 4461
rect 126 4432 129 4458
rect 155 4432 158 4458
rect 126 4429 158 4432
rect 135 4385 150 4429
rect 128 4382 154 4385
rect 128 4353 154 4356
rect 135 4248 150 4353
rect 127 4245 159 4248
rect 127 4219 130 4245
rect 156 4219 159 4245
rect 127 4216 159 4219
rect 135 4162 150 4216
rect 127 4159 159 4162
rect 127 4133 130 4159
rect 156 4133 159 4159
rect 127 4130 159 4133
rect 135 4088 150 4130
rect 128 4085 154 4088
rect 128 4056 154 4059
rect 135 4005 150 4056
rect 127 4002 159 4005
rect 127 3976 130 4002
rect 156 3976 159 4002
rect 127 3973 159 3976
rect 135 3921 150 3973
rect 127 3918 159 3921
rect 127 3892 130 3918
rect 156 3892 159 3918
rect 127 3889 159 3892
rect 135 3847 150 3889
rect 129 3844 155 3847
rect 129 3815 155 3818
rect 135 3606 150 3815
rect 129 3603 155 3606
rect 129 3574 155 3577
rect 135 3365 150 3574
rect 129 3362 155 3365
rect 129 3333 155 3336
rect 135 3124 150 3333
rect 129 3121 155 3124
rect 129 3092 155 3095
rect 135 2883 150 3092
rect 129 2880 155 2883
rect 129 2851 155 2854
rect 135 2602 150 2851
rect 128 2599 154 2602
rect 128 2570 154 2573
rect 135 2361 150 2570
rect 129 2358 155 2361
rect 129 2329 155 2332
rect 135 2120 150 2329
rect 129 2117 155 2120
rect 129 2088 155 2091
rect 135 1879 150 2088
rect 129 1876 155 1879
rect 129 1847 155 1850
rect 135 1638 150 1847
rect 129 1635 155 1638
rect 129 1606 155 1609
rect 135 1397 150 1606
rect 129 1394 155 1397
rect 129 1365 155 1368
rect 135 1156 150 1365
rect 128 1153 154 1156
rect 128 1124 154 1127
rect 135 915 150 1124
rect 129 912 155 915
rect 129 883 155 886
rect 135 633 150 883
rect 128 630 154 633
rect 128 601 154 604
rect 135 392 150 601
rect 130 389 156 392
rect 130 360 156 363
rect 135 151 150 360
rect 129 148 155 151
rect 129 119 155 122
rect 135 -90 150 119
rect 126 -93 158 -90
rect 126 -119 129 -93
rect 155 -119 158 -93
rect 126 -122 158 -119
rect 135 -175 150 -122
rect 126 -178 158 -175
rect 126 -204 129 -178
rect 155 -204 158 -178
rect 126 -207 158 -204
rect 135 -254 150 -207
rect 126 -257 158 -254
rect 126 -283 129 -257
rect 155 -283 158 -257
rect 126 -286 158 -283
rect 135 -334 150 -286
rect 126 -360 129 -334
rect 155 -360 158 -334
rect 135 -413 150 -360
rect 126 -416 158 -413
rect 126 -442 129 -416
rect 155 -442 158 -416
rect 126 -445 158 -442
rect 135 -492 150 -445
rect 127 -495 159 -492
rect 127 -521 130 -495
rect 156 -521 159 -495
rect 127 -524 159 -521
rect 135 -572 150 -524
rect 129 -575 155 -572
rect 129 -604 155 -601
rect 135 -715 150 -604
rect 126 -718 158 -715
rect 126 -744 129 -718
rect 155 -744 158 -718
rect 126 -747 158 -744
rect 135 -795 150 -747
rect 126 -798 158 -795
rect 126 -824 129 -798
rect 155 -824 158 -798
rect 126 -827 158 -824
rect 135 -872 150 -827
rect 126 -875 158 -872
rect 126 -901 129 -875
rect 155 -901 158 -875
rect 126 -904 158 -901
rect 135 -952 150 -904
rect 126 -955 158 -952
rect 126 -981 129 -955
rect 155 -981 158 -955
rect 126 -984 158 -981
rect 135 -1039 150 -984
rect 127 -1042 159 -1039
rect 127 -1068 130 -1042
rect 156 -1068 159 -1042
rect 127 -1071 159 -1068
rect 135 -1113 150 -1071
rect 129 -1116 155 -1113
rect 129 -1145 155 -1142
rect 135 -1890 150 -1145
rect 129 -1893 155 -1890
rect 129 -1922 155 -1919
rect -4180 -2034 -4150 -2029
rect -4180 -2069 -4150 -2064
rect -40 -2030 0 -2025
rect 135 -2030 150 -1922
rect -40 -2060 -35 -2030
rect -5 -2060 0 -2030
rect -40 -2065 0 -2060
rect 126 -2033 159 -2030
rect 126 -2059 130 -2033
rect 156 -2059 159 -2033
rect 126 -2062 159 -2059
rect -4314 -3063 -4284 -3058
rect -4314 -3098 -4284 -3093
rect -4172 -4343 -4158 -2069
rect 234 -2098 248 5356
rect 519 5069 559 5074
rect 519 5039 524 5069
rect 554 5039 559 5069
rect 519 5034 559 5039
rect 596 -607 626 -602
rect 596 -642 626 -637
rect 602 -1383 619 -642
rect 594 -1386 626 -1383
rect 594 -1412 597 -1386
rect 623 -1412 626 -1386
rect 594 -1415 626 -1412
rect 815 -2096 829 5345
rect 1095 5069 1135 5074
rect 1095 5039 1100 5069
rect 1130 5039 1135 5069
rect 1095 5034 1135 5039
rect 1171 -734 1201 -729
rect 1171 -769 1201 -764
rect 1177 -1384 1194 -769
rect 1169 -1387 1201 -1384
rect 1169 -1413 1172 -1387
rect 1198 -1413 1201 -1387
rect 1169 -1416 1201 -1413
rect 225 -2101 257 -2098
rect 225 -2127 228 -2101
rect 254 -2127 257 -2101
rect 225 -2130 257 -2127
rect 806 -2099 838 -2096
rect 1386 -2097 1400 5341
rect 1670 5069 1710 5074
rect 1670 5039 1675 5069
rect 1705 5039 1710 5069
rect 1670 5034 1710 5039
rect 1751 -871 1781 -866
rect 1751 -906 1781 -901
rect 1752 -1386 1769 -906
rect 1744 -1389 1776 -1386
rect 1744 -1415 1747 -1389
rect 1773 -1415 1776 -1389
rect 1744 -1418 1776 -1415
rect 806 -2125 809 -2099
rect 835 -2125 838 -2099
rect 806 -2128 838 -2125
rect 1378 -2100 1410 -2097
rect 1964 -2099 1978 5342
rect 2243 5069 2283 5074
rect 2243 5039 2248 5069
rect 2278 5039 2283 5069
rect 2243 5034 2283 5039
rect 2321 -988 2351 -983
rect 2321 -1023 2351 -1018
rect 2327 -1386 2344 -1023
rect 2319 -1389 2351 -1386
rect 2319 -1415 2322 -1389
rect 2348 -1415 2351 -1389
rect 2319 -1418 2351 -1415
rect 2537 -2099 2551 5342
rect 2819 5069 2859 5074
rect 2819 5039 2824 5069
rect 2854 5039 2859 5069
rect 2819 5034 2859 5039
rect 2896 -1113 2926 -1108
rect 2896 -1148 2926 -1143
rect 2902 -1384 2919 -1148
rect 2894 -1387 2926 -1384
rect 2894 -1413 2897 -1387
rect 2923 -1413 2926 -1387
rect 2894 -1416 2926 -1413
rect 1378 -2126 1381 -2100
rect 1407 -2126 1410 -2100
rect 1378 -2129 1410 -2126
rect 1956 -2102 1988 -2099
rect 1956 -2128 1959 -2102
rect 1985 -2128 1988 -2102
rect 1956 -2131 1988 -2128
rect 2531 -2102 2563 -2099
rect 3110 -2101 3124 5340
rect 3393 5069 3433 5074
rect 3393 5039 3398 5069
rect 3428 5039 3433 5069
rect 3393 5034 3433 5039
rect 3471 -1258 3501 -1253
rect 3471 -1293 3501 -1288
rect 3477 -1381 3494 -1293
rect 3469 -1384 3501 -1381
rect 3469 -1410 3472 -1384
rect 3498 -1410 3501 -1384
rect 3469 -1413 3501 -1410
rect 3686 -2100 3700 5341
rect 3968 5069 4008 5074
rect 3968 5039 3973 5069
rect 4003 5039 4008 5069
rect 3968 5034 4008 5039
rect 4040 -1380 4080 -1375
rect 4040 -1410 4045 -1380
rect 4075 -1410 4080 -1380
rect 4040 -1415 4080 -1410
rect 4264 -2099 4278 5342
rect 4543 5069 4583 5074
rect 4543 5039 4548 5069
rect 4578 5039 4583 5069
rect 4543 5034 4583 5039
rect 4619 -1382 4651 -1379
rect 4619 -1408 4622 -1382
rect 4648 -1408 4651 -1382
rect 4619 -1411 4651 -1408
rect 4627 -1463 4644 -1411
rect 4621 -1468 4651 -1463
rect 4621 -1503 4651 -1498
rect 4837 -2098 4851 5342
rect 5118 5069 5158 5074
rect 5118 5039 5123 5069
rect 5153 5039 5158 5069
rect 5118 5034 5158 5039
rect 5194 -1387 5226 -1384
rect 5194 -1413 5197 -1387
rect 5223 -1413 5226 -1387
rect 5194 -1416 5226 -1413
rect 5202 -1546 5219 -1416
rect 5196 -1551 5226 -1546
rect 5196 -1586 5226 -1581
rect 2531 -2128 2534 -2102
rect 2560 -2128 2563 -2102
rect 2531 -2131 2563 -2128
rect 3102 -2104 3134 -2101
rect 3102 -2130 3105 -2104
rect 3131 -2130 3134 -2104
rect 3102 -2133 3134 -2130
rect 3679 -2103 3711 -2100
rect 3679 -2129 3682 -2103
rect 3708 -2129 3711 -2103
rect 3679 -2132 3711 -2129
rect 4259 -2102 4291 -2099
rect 4259 -2128 4262 -2102
rect 4288 -2128 4291 -2102
rect 4259 -2131 4291 -2128
rect 4829 -2101 4861 -2098
rect 5412 -2100 5426 5340
rect 5694 5069 5734 5074
rect 5694 5039 5699 5069
rect 5729 5039 5734 5069
rect 5694 5034 5734 5039
rect 5769 -1384 5801 -1381
rect 5769 -1410 5772 -1384
rect 5798 -1410 5801 -1384
rect 5769 -1413 5801 -1410
rect 5777 -1624 5794 -1413
rect 5771 -1629 5801 -1624
rect 5771 -1664 5801 -1659
rect 5988 -2098 6002 5341
rect 6269 5068 6309 5073
rect 6269 5038 6274 5068
rect 6304 5038 6309 5068
rect 6269 5033 6309 5038
rect 6344 -1388 6376 -1385
rect 6344 -1414 6347 -1388
rect 6373 -1414 6376 -1388
rect 6344 -1417 6376 -1414
rect 6352 -1710 6369 -1417
rect 6346 -1715 6376 -1710
rect 6346 -1750 6376 -1745
rect 4829 -2127 4832 -2101
rect 4858 -2127 4861 -2101
rect 4829 -2130 4861 -2127
rect 5406 -2103 5438 -2100
rect 5406 -2129 5409 -2103
rect 5435 -2129 5438 -2103
rect 5406 -2132 5438 -2129
rect 5980 -2101 6012 -2098
rect 6561 -2099 6575 5341
rect 6843 5069 6883 5074
rect 6843 5039 6848 5069
rect 6878 5039 6883 5069
rect 6843 5034 6883 5039
rect 6919 -1389 6951 -1386
rect 6919 -1415 6922 -1389
rect 6948 -1415 6951 -1389
rect 6919 -1418 6951 -1415
rect 6927 -1790 6944 -1418
rect 6921 -1795 6951 -1790
rect 6921 -1830 6951 -1825
rect 5980 -2127 5983 -2101
rect 6009 -2127 6012 -2101
rect 5980 -2130 6012 -2127
rect 6553 -2102 6585 -2099
rect 7136 -2100 7150 5341
rect 7418 5069 7458 5074
rect 7418 5039 7423 5069
rect 7453 5039 7458 5069
rect 7418 5034 7458 5039
rect 7494 -1385 7526 -1382
rect 7494 -1411 7497 -1385
rect 7523 -1411 7526 -1385
rect 7494 -1414 7526 -1411
rect 7502 -1870 7519 -1414
rect 7496 -1875 7526 -1870
rect 7496 -1910 7526 -1905
rect 7711 -2100 7725 5342
rect 7993 5069 8033 5074
rect 7993 5039 7998 5069
rect 8028 5039 8033 5069
rect 7993 5034 8033 5039
rect 8069 -1389 8101 -1386
rect 8069 -1415 8072 -1389
rect 8098 -1415 8101 -1389
rect 8069 -1418 8101 -1415
rect 8077 -1935 8094 -1418
rect 8071 -1940 8101 -1935
rect 8071 -1975 8101 -1970
rect 6553 -2128 6556 -2102
rect 6582 -2128 6585 -2102
rect 6553 -2131 6585 -2128
rect 7130 -2103 7162 -2100
rect 7130 -2129 7133 -2103
rect 7159 -2129 7162 -2103
rect 7130 -2132 7162 -2129
rect 7706 -2103 7738 -2100
rect 8288 -2102 8302 5342
rect 8567 5069 8607 5074
rect 8567 5039 8572 5069
rect 8602 5039 8607 5069
rect 8567 5034 8607 5039
rect 8644 -1385 8676 -1382
rect 8644 -1411 8647 -1385
rect 8673 -1411 8676 -1385
rect 8644 -1414 8676 -1411
rect 8652 -2049 8669 -1414
rect 8646 -2054 8676 -2049
rect 8646 -2089 8676 -2084
rect 8863 -2102 8877 5342
rect 9142 5069 9182 5074
rect 9142 5039 9147 5069
rect 9177 5039 9182 5069
rect 9142 5034 9182 5039
rect 9219 -1386 9251 -1383
rect 9219 -1412 9222 -1386
rect 9248 -1412 9251 -1386
rect 9219 -1415 9251 -1412
rect 7706 -2129 7709 -2103
rect 7735 -2129 7738 -2103
rect 7706 -2132 7738 -2129
rect 8279 -2105 8311 -2102
rect 8279 -2131 8282 -2105
rect 8308 -2131 8311 -2105
rect 8279 -2134 8311 -2131
rect 8854 -2105 8886 -2102
rect 8854 -2131 8857 -2105
rect 8883 -2131 8886 -2105
rect 8854 -2134 8886 -2131
rect 9227 -2138 9244 -1415
rect 9221 -2143 9251 -2138
rect 9221 -2178 9251 -2173
rect 305 -2271 319 -2242
rect 296 -2274 328 -2271
rect 296 -2300 299 -2274
rect 325 -2300 328 -2274
rect 296 -2303 328 -2300
rect 532 -2338 546 -2242
rect 758 -2271 772 -2255
rect 880 -2271 894 -2256
rect 749 -2274 781 -2271
rect 749 -2300 752 -2274
rect 778 -2300 781 -2274
rect 749 -2303 781 -2300
rect 871 -2274 903 -2271
rect 871 -2300 874 -2274
rect 900 -2300 903 -2274
rect 871 -2303 903 -2300
rect 806 -2320 846 -2315
rect 523 -2341 555 -2338
rect 523 -2367 526 -2341
rect 552 -2367 555 -2341
rect 806 -2350 811 -2320
rect 841 -2350 846 -2320
rect 1107 -2339 1121 -2242
rect 1333 -2271 1347 -2256
rect 1455 -2271 1469 -2256
rect 1324 -2274 1356 -2271
rect 1324 -2300 1327 -2274
rect 1353 -2300 1356 -2274
rect 1324 -2303 1356 -2300
rect 1446 -2274 1478 -2271
rect 1446 -2300 1449 -2274
rect 1475 -2300 1478 -2274
rect 1446 -2303 1478 -2300
rect 806 -2355 846 -2350
rect 1098 -2342 1130 -2339
rect 523 -2370 555 -2367
rect 1098 -2368 1101 -2342
rect 1127 -2368 1130 -2342
rect 1682 -2344 1696 -2256
rect 1908 -2271 1922 -2256
rect 2030 -2271 2044 -2256
rect 1899 -2274 1931 -2271
rect 1899 -2300 1902 -2274
rect 1928 -2300 1931 -2274
rect 1899 -2303 1931 -2300
rect 2021 -2274 2053 -2271
rect 2021 -2300 2024 -2274
rect 2050 -2300 2053 -2274
rect 2021 -2303 2053 -2300
rect 1955 -2321 1995 -2316
rect 1098 -2371 1130 -2368
rect 1673 -2347 1705 -2344
rect 1673 -2373 1676 -2347
rect 1702 -2373 1705 -2347
rect 1955 -2351 1960 -2321
rect 1990 -2351 1995 -2321
rect 2257 -2344 2271 -2256
rect 2483 -2271 2497 -2256
rect 2605 -2271 2619 -2256
rect 2474 -2274 2506 -2271
rect 2474 -2300 2477 -2274
rect 2503 -2300 2506 -2274
rect 2474 -2303 2506 -2300
rect 2596 -2274 2628 -2271
rect 2596 -2300 2599 -2274
rect 2625 -2300 2628 -2274
rect 2596 -2303 2628 -2300
rect 2832 -2344 2846 -2256
rect 3058 -2271 3072 -2256
rect 3180 -2271 3194 -2256
rect 3049 -2274 3081 -2271
rect 3049 -2300 3052 -2274
rect 3078 -2300 3081 -2274
rect 3049 -2303 3081 -2300
rect 3171 -2274 3203 -2271
rect 3171 -2300 3174 -2274
rect 3200 -2300 3203 -2274
rect 3171 -2303 3203 -2300
rect 3098 -2322 3138 -2317
rect 1955 -2356 1995 -2351
rect 2248 -2347 2280 -2344
rect 1673 -2376 1705 -2373
rect 2248 -2373 2251 -2347
rect 2277 -2373 2280 -2347
rect 2248 -2376 2280 -2373
rect 2823 -2347 2855 -2344
rect 2823 -2373 2826 -2347
rect 2852 -2373 2855 -2347
rect 3098 -2352 3103 -2322
rect 3133 -2352 3138 -2322
rect 3407 -2344 3421 -2256
rect 3633 -2271 3647 -2256
rect 3755 -2271 3769 -2256
rect 3624 -2274 3656 -2271
rect 3624 -2300 3627 -2274
rect 3653 -2300 3656 -2274
rect 3624 -2303 3656 -2300
rect 3746 -2274 3778 -2271
rect 3746 -2300 3749 -2274
rect 3775 -2300 3778 -2274
rect 3746 -2303 3778 -2300
rect 3982 -2344 3996 -2256
rect 4208 -2271 4222 -2256
rect 4330 -2271 4344 -2256
rect 4199 -2274 4231 -2271
rect 4199 -2300 4202 -2274
rect 4228 -2300 4231 -2274
rect 4199 -2303 4231 -2300
rect 4321 -2274 4353 -2271
rect 4321 -2300 4324 -2274
rect 4350 -2300 4353 -2274
rect 4321 -2303 4353 -2300
rect 4255 -2323 4295 -2318
rect 3098 -2357 3138 -2352
rect 3398 -2347 3430 -2344
rect 2823 -2376 2855 -2373
rect 3398 -2373 3401 -2347
rect 3427 -2373 3430 -2347
rect 3398 -2376 3430 -2373
rect 3973 -2347 4005 -2344
rect 3973 -2373 3976 -2347
rect 4002 -2373 4005 -2347
rect 4255 -2353 4260 -2323
rect 4290 -2353 4295 -2323
rect 4557 -2344 4571 -2256
rect 4783 -2271 4797 -2256
rect 4905 -2271 4919 -2256
rect 4774 -2274 4806 -2271
rect 4774 -2300 4777 -2274
rect 4803 -2300 4806 -2274
rect 4774 -2303 4806 -2300
rect 4896 -2274 4928 -2271
rect 4896 -2300 4899 -2274
rect 4925 -2300 4928 -2274
rect 4896 -2303 4928 -2300
rect 5132 -2344 5146 -2256
rect 5358 -2271 5372 -2256
rect 5480 -2271 5494 -2256
rect 5349 -2274 5381 -2271
rect 5349 -2300 5352 -2274
rect 5378 -2300 5381 -2274
rect 5349 -2303 5381 -2300
rect 5471 -2274 5503 -2271
rect 5471 -2300 5474 -2274
rect 5500 -2300 5503 -2274
rect 5471 -2303 5503 -2300
rect 5395 -2321 5435 -2316
rect 4255 -2358 4295 -2353
rect 4548 -2347 4580 -2344
rect 3973 -2376 4005 -2373
rect 4548 -2373 4551 -2347
rect 4577 -2373 4580 -2347
rect 4548 -2376 4580 -2373
rect 5123 -2347 5155 -2344
rect 5123 -2373 5126 -2347
rect 5152 -2373 5155 -2347
rect 5395 -2351 5400 -2321
rect 5430 -2351 5435 -2321
rect 5707 -2344 5721 -2256
rect 5933 -2271 5947 -2256
rect 6055 -2271 6069 -2256
rect 5924 -2274 5956 -2271
rect 5924 -2300 5927 -2274
rect 5953 -2300 5956 -2274
rect 5924 -2303 5956 -2300
rect 6046 -2274 6078 -2271
rect 6046 -2300 6049 -2274
rect 6075 -2300 6078 -2274
rect 6046 -2303 6078 -2300
rect 6282 -2344 6296 -2256
rect 6508 -2271 6522 -2256
rect 6630 -2271 6644 -2256
rect 6499 -2274 6531 -2271
rect 6499 -2300 6502 -2274
rect 6528 -2300 6531 -2274
rect 6499 -2303 6531 -2300
rect 6621 -2274 6653 -2271
rect 6621 -2300 6624 -2274
rect 6650 -2300 6653 -2274
rect 6621 -2303 6653 -2300
rect 6563 -2321 6603 -2316
rect 5395 -2356 5435 -2351
rect 5698 -2347 5730 -2344
rect 5123 -2376 5155 -2373
rect 5698 -2373 5701 -2347
rect 5727 -2373 5730 -2347
rect 5698 -2376 5730 -2373
rect 6273 -2347 6305 -2344
rect 6273 -2373 6276 -2347
rect 6302 -2373 6305 -2347
rect 6563 -2351 6568 -2321
rect 6598 -2351 6603 -2321
rect 6857 -2344 6871 -2256
rect 7083 -2271 7097 -2256
rect 7205 -2271 7219 -2256
rect 7074 -2274 7106 -2271
rect 7074 -2300 7077 -2274
rect 7103 -2300 7106 -2274
rect 7074 -2303 7106 -2300
rect 7196 -2274 7228 -2271
rect 7196 -2300 7199 -2274
rect 7225 -2300 7228 -2274
rect 7196 -2303 7228 -2300
rect 7432 -2344 7446 -2256
rect 7658 -2271 7672 -2256
rect 7780 -2271 7794 -2256
rect 7649 -2274 7681 -2271
rect 7649 -2300 7652 -2274
rect 7678 -2300 7681 -2274
rect 7649 -2303 7681 -2300
rect 7771 -2274 7803 -2271
rect 7771 -2300 7774 -2274
rect 7800 -2300 7803 -2274
rect 7771 -2303 7803 -2300
rect 7708 -2321 7748 -2316
rect 6563 -2356 6603 -2351
rect 6848 -2347 6880 -2344
rect 6273 -2376 6305 -2373
rect 6848 -2373 6851 -2347
rect 6877 -2373 6880 -2347
rect 6848 -2376 6880 -2373
rect 7423 -2347 7455 -2344
rect 7423 -2373 7426 -2347
rect 7452 -2373 7455 -2347
rect 7708 -2351 7713 -2321
rect 7743 -2351 7748 -2321
rect 8007 -2344 8021 -2256
rect 8233 -2271 8247 -2256
rect 8355 -2271 8369 -2256
rect 8224 -2274 8256 -2271
rect 8224 -2300 8227 -2274
rect 8253 -2300 8256 -2274
rect 8224 -2303 8256 -2300
rect 8346 -2274 8378 -2271
rect 8346 -2300 8349 -2274
rect 8375 -2300 8378 -2274
rect 8346 -2303 8378 -2300
rect 8582 -2344 8596 -2256
rect 8808 -2271 8822 -2256
rect 8930 -2271 8944 -2256
rect 8799 -2274 8831 -2271
rect 8799 -2300 8802 -2274
rect 8828 -2300 8831 -2274
rect 8799 -2303 8831 -2300
rect 8921 -2274 8953 -2271
rect 8921 -2300 8924 -2274
rect 8950 -2300 8953 -2274
rect 8921 -2303 8953 -2300
rect 8865 -2319 8905 -2314
rect 7708 -2356 7748 -2351
rect 7998 -2347 8030 -2344
rect 7423 -2376 7455 -2373
rect 7998 -2373 8001 -2347
rect 8027 -2373 8030 -2347
rect 7998 -2376 8030 -2373
rect 8573 -2347 8605 -2344
rect 8573 -2373 8576 -2347
rect 8602 -2373 8605 -2347
rect 8865 -2349 8870 -2319
rect 8900 -2349 8905 -2319
rect 9157 -2344 9171 -2256
rect 9383 -2271 9397 -2256
rect 9374 -2274 9406 -2271
rect 9374 -2300 9377 -2274
rect 9403 -2300 9406 -2274
rect 9374 -2303 9406 -2300
rect 8865 -2354 8905 -2349
rect 9148 -2347 9180 -2344
rect 8573 -2376 8605 -2373
rect 9148 -2373 9151 -2347
rect 9177 -2373 9180 -2347
rect 9148 -2376 9180 -2373
rect 730 -2419 770 -2414
rect 730 -2449 735 -2419
rect 765 -2449 770 -2419
rect 730 -2454 770 -2449
rect 885 -2419 925 -2414
rect 885 -2449 890 -2419
rect 920 -2449 925 -2419
rect 885 -2454 925 -2449
rect 1880 -2419 1920 -2414
rect 1880 -2449 1885 -2419
rect 1915 -2449 1920 -2419
rect 1880 -2454 1920 -2449
rect 2035 -2419 2075 -2414
rect 2035 -2449 2040 -2419
rect 2070 -2449 2075 -2419
rect 2035 -2454 2075 -2449
rect 3030 -2419 3070 -2414
rect 3030 -2449 3035 -2419
rect 3065 -2449 3070 -2419
rect 3030 -2454 3070 -2449
rect 3184 -2419 3224 -2414
rect 3184 -2449 3189 -2419
rect 3219 -2449 3224 -2419
rect 3184 -2454 3224 -2449
rect 4177 -2419 4217 -2414
rect 4177 -2449 4182 -2419
rect 4212 -2449 4217 -2419
rect 4177 -2454 4217 -2449
rect 4336 -2420 4376 -2415
rect 4336 -2450 4341 -2420
rect 4371 -2450 4376 -2420
rect 4336 -2455 4376 -2450
rect 5329 -2419 5369 -2414
rect 5329 -2449 5334 -2419
rect 5364 -2449 5369 -2419
rect 5329 -2454 5369 -2449
rect 5484 -2419 5524 -2414
rect 5484 -2449 5489 -2419
rect 5519 -2449 5524 -2419
rect 5484 -2454 5524 -2449
rect 6480 -2420 6520 -2415
rect 6480 -2450 6485 -2420
rect 6515 -2450 6520 -2420
rect 6480 -2455 6520 -2450
rect 6633 -2420 6673 -2415
rect 6633 -2450 6638 -2420
rect 6668 -2450 6673 -2420
rect 6633 -2455 6673 -2450
rect 7631 -2419 7671 -2414
rect 7631 -2449 7636 -2419
rect 7666 -2449 7671 -2419
rect 7631 -2454 7671 -2449
rect 7784 -2419 7824 -2414
rect 7784 -2449 7789 -2419
rect 7819 -2449 7824 -2419
rect 7784 -2454 7824 -2449
rect 8780 -2418 8820 -2414
rect 8780 -2448 8785 -2418
rect 8815 -2448 8820 -2418
rect 8780 -2454 8820 -2448
rect 8932 -2419 8972 -2413
rect 8932 -2449 8937 -2419
rect 8967 -2449 8972 -2419
rect 8932 -2454 8972 -2449
rect -3927 -2458 -3895 -2455
rect -3927 -2484 -3924 -2458
rect -3898 -2484 -3895 -2458
rect -3927 -2487 -3895 -2484
rect -3988 -3125 -3962 -3122
rect -3988 -3154 -3962 -3151
rect -4054 -3628 -4028 -3625
rect -4054 -3657 -4028 -3654
rect -4120 -3668 -4094 -3665
rect -4120 -3697 -4094 -3694
rect -4178 -4346 -4152 -4343
rect -4178 -4375 -4152 -4372
rect -4114 -5311 -4100 -3697
rect -4123 -5314 -4091 -5311
rect -4123 -5340 -4120 -5314
rect -4094 -5340 -4091 -5314
rect -4123 -5343 -4091 -5340
rect -4114 -6398 -4100 -5343
rect -4048 -5351 -4034 -3657
rect -4054 -5354 -4028 -5351
rect -4054 -5383 -4028 -5380
rect -4048 -6358 -4034 -5383
rect -3982 -5854 -3968 -3154
rect -3918 -4128 -3904 -2487
rect 1154 -2489 1194 -2484
rect 461 -2496 501 -2491
rect 461 -2526 466 -2496
rect 496 -2526 501 -2496
rect 1154 -2519 1159 -2489
rect 1189 -2519 1194 -2489
rect 1154 -2524 1194 -2519
rect 1610 -2488 1650 -2483
rect 1610 -2518 1615 -2488
rect 1645 -2518 1650 -2488
rect 1610 -2523 1650 -2518
rect 2303 -2493 2343 -2488
rect 2303 -2523 2308 -2493
rect 2338 -2523 2343 -2493
rect 461 -2531 501 -2526
rect 2303 -2528 2343 -2523
rect 2762 -2494 2802 -2489
rect 2762 -2524 2767 -2494
rect 2797 -2524 2802 -2494
rect 2762 -2529 2802 -2524
rect 3454 -2492 3494 -2487
rect 3454 -2522 3459 -2492
rect 3489 -2522 3494 -2492
rect 3454 -2527 3494 -2522
rect 3912 -2494 3952 -2489
rect 5061 -2490 5101 -2485
rect 3912 -2524 3917 -2494
rect 3947 -2524 3952 -2494
rect 3912 -2529 3952 -2524
rect 4603 -2496 4643 -2491
rect 4603 -2526 4608 -2496
rect 4638 -2526 4643 -2496
rect 5061 -2520 5066 -2490
rect 5096 -2520 5101 -2490
rect 5061 -2525 5101 -2520
rect 5754 -2492 5794 -2487
rect 5754 -2522 5759 -2492
rect 5789 -2522 5794 -2492
rect 4603 -2531 4643 -2526
rect 5754 -2527 5794 -2522
rect 6211 -2488 6251 -2483
rect 6211 -2518 6216 -2488
rect 6246 -2518 6251 -2488
rect 6211 -2523 6251 -2518
rect 6903 -2492 6943 -2487
rect 6903 -2522 6908 -2492
rect 6938 -2522 6943 -2492
rect 6903 -2527 6943 -2522
rect 7361 -2492 7401 -2487
rect 7361 -2522 7366 -2492
rect 7396 -2522 7401 -2492
rect 7361 -2527 7401 -2522
rect 8053 -2495 8093 -2490
rect 8053 -2525 8058 -2495
rect 8088 -2525 8093 -2495
rect 8053 -2530 8093 -2525
rect 8511 -2493 8551 -2489
rect 8511 -2523 8516 -2493
rect 8546 -2523 8551 -2493
rect 8511 -2529 8551 -2523
rect 9203 -2491 9239 -2487
rect 9203 -2521 9206 -2491
rect 9236 -2521 9239 -2491
rect 9203 -2525 9239 -2521
rect 13532 -2537 13558 -2534
rect -2747 -2540 -2715 -2537
rect -2747 -2566 -2744 -2540
rect -2718 -2566 -2715 -2540
rect 13532 -2566 13558 -2563
rect -2747 -2569 -2715 -2566
rect -3524 -3067 -3494 -3062
rect -3524 -3102 -3494 -3097
rect -3516 -3134 -3502 -3102
rect -3148 -3584 -3122 -3581
rect -3148 -3613 -3122 -3610
rect -3930 -4131 -3892 -4128
rect -3930 -4163 -3927 -4131
rect -3895 -4163 -3892 -4131
rect -3930 -4166 -3892 -4163
rect -3913 -4346 -3887 -4343
rect -3913 -4375 -3887 -4372
rect -3907 -4633 -3893 -4375
rect -3913 -4636 -3887 -4633
rect -3913 -4665 -3887 -4662
rect -3987 -5857 -3961 -5854
rect -3987 -5886 -3961 -5883
rect -4057 -6361 -4025 -6358
rect -4057 -6387 -4054 -6361
rect -4028 -6387 -4025 -6361
rect -4057 -6390 -4025 -6387
rect -4123 -6401 -4091 -6398
rect -4123 -6427 -4120 -6401
rect -4094 -6427 -4091 -6401
rect -4123 -6430 -4091 -6427
rect -4114 -8044 -4100 -6430
rect -4123 -8047 -4091 -8044
rect -4123 -8073 -4120 -8047
rect -4094 -8073 -4091 -8047
rect -4123 -8076 -4091 -8073
rect -4114 -9025 -4100 -8076
rect -4048 -8084 -4034 -6390
rect -4057 -8087 -4025 -8084
rect -4057 -8113 -4054 -8087
rect -4028 -8113 -4025 -8087
rect -4057 -8116 -4025 -8113
rect -4048 -9025 -4034 -8116
rect -3982 -8587 -3968 -5886
rect -3907 -7076 -3893 -4665
rect -3913 -7079 -3887 -7076
rect -3913 -7108 -3887 -7105
rect -3907 -7369 -3893 -7108
rect -3916 -7395 -3913 -7369
rect -3887 -7395 -3884 -7369
rect -3991 -8590 -3959 -8587
rect -3991 -8616 -3988 -8590
rect -3962 -8616 -3959 -8590
rect -3991 -8619 -3959 -8616
rect -3982 -9025 -3968 -8619
rect -3142 -9017 -3128 -3613
rect -2739 -4132 -2722 -2569
rect -1565 -2603 -1539 -2600
rect 12583 -2613 12586 -2587
rect 12612 -2613 12615 -2587
rect -1565 -2632 -1539 -2629
rect -2374 -3067 -2344 -3062
rect -2374 -3102 -2344 -3097
rect -2366 -3131 -2352 -3102
rect -1993 -3584 -1967 -3581
rect -1993 -3613 -1967 -3610
rect -2746 -4135 -2714 -4132
rect -2746 -4161 -2743 -4135
rect -2717 -4161 -2714 -4135
rect -2746 -4164 -2714 -4161
rect -3107 -5397 -3081 -5394
rect -3107 -5426 -3081 -5423
rect -3101 -9017 -3087 -5426
rect -3067 -6317 -3041 -6314
rect -3067 -6346 -3041 -6343
rect -3061 -9017 -3047 -6346
rect -3026 -8130 -3000 -8127
rect -3026 -8159 -3000 -8156
rect -3020 -9017 -3006 -8159
rect -1987 -9009 -1973 -3613
rect -1560 -4132 -1543 -2632
rect 11420 -2663 11423 -2637
rect 11449 -2663 11452 -2637
rect -387 -2678 -361 -2675
rect -387 -2707 -361 -2704
rect -1192 -3066 -1162 -3061
rect -1192 -3101 -1162 -3096
rect -1184 -3131 -1170 -3101
rect -824 -3584 -798 -3581
rect -824 -3613 -798 -3610
rect -1564 -4135 -1538 -4132
rect -1564 -4164 -1538 -4161
rect -1953 -5397 -1927 -5394
rect -1953 -5426 -1927 -5423
rect -1947 -9009 -1933 -5426
rect -1914 -6317 -1882 -6314
rect -1914 -6343 -1911 -6317
rect -1885 -6343 -1882 -6317
rect -1914 -6346 -1882 -6343
rect -1905 -9009 -1891 -6346
rect -1870 -8130 -1844 -8127
rect -1870 -8159 -1844 -8156
rect -1864 -9009 -1850 -8159
rect -818 -8986 -804 -3613
rect -382 -4132 -365 -2707
rect 10207 -2726 10210 -2700
rect 10236 -2726 10239 -2700
rect 808 -2749 840 -2746
rect 808 -2775 811 -2749
rect 837 -2775 840 -2749
rect 808 -2778 840 -2775
rect -11 -3071 19 -3066
rect -11 -3106 19 -3101
rect -3 -3131 11 -3106
rect 367 -3584 393 -3581
rect 367 -3613 393 -3610
rect -386 -4135 -360 -4132
rect -386 -4164 -360 -4161
rect -784 -5397 -758 -5394
rect -784 -5426 -758 -5423
rect -778 -8986 -764 -5426
rect -745 -6317 -713 -6314
rect -745 -6343 -742 -6317
rect -716 -6343 -713 -6317
rect -745 -6346 -713 -6343
rect -736 -8986 -722 -6346
rect -701 -8130 -675 -8127
rect -701 -8159 -675 -8156
rect -695 -8986 -681 -8159
rect 373 -8978 387 -3613
rect 816 -4132 833 -2778
rect 9033 -2789 9036 -2763
rect 9062 -2789 9065 -2763
rect 1975 -2829 2007 -2826
rect 1975 -2855 1978 -2829
rect 2004 -2855 2007 -2829
rect 1975 -2858 2007 -2855
rect 7848 -2835 7874 -2832
rect 1170 -3069 1200 -3064
rect 1170 -3104 1200 -3099
rect 1178 -3132 1192 -3104
rect 1544 -3584 1570 -3581
rect 1544 -3613 1570 -3610
rect 809 -4135 841 -4132
rect 809 -4161 812 -4135
rect 838 -4161 841 -4135
rect 809 -4164 841 -4161
rect 407 -5397 433 -5394
rect 407 -5426 433 -5423
rect 413 -8978 427 -5426
rect 446 -6317 478 -6314
rect 446 -6343 449 -6317
rect 475 -6343 478 -6317
rect 446 -6346 478 -6343
rect 455 -8978 469 -6346
rect 490 -8130 516 -8127
rect 490 -8159 516 -8156
rect 496 -8978 510 -8159
rect 1550 -8995 1564 -3613
rect 1983 -4131 2000 -2858
rect 7848 -2864 7874 -2861
rect 3134 -2913 3166 -2910
rect 3134 -2939 3137 -2913
rect 3163 -2939 3166 -2913
rect 3134 -2942 3166 -2939
rect 6646 -2915 6672 -2912
rect 2352 -3070 2382 -3065
rect 2352 -3105 2382 -3100
rect 2360 -3131 2374 -3105
rect 2721 -3584 2747 -3581
rect 2721 -3613 2747 -3610
rect 1975 -4134 2008 -4131
rect 1975 -4160 1979 -4134
rect 2005 -4160 2008 -4134
rect 1975 -4163 2008 -4160
rect 1584 -5397 1610 -5394
rect 1584 -5426 1610 -5423
rect 1590 -8995 1604 -5426
rect 1623 -6317 1655 -6314
rect 1623 -6343 1626 -6317
rect 1652 -6343 1655 -6317
rect 1623 -6346 1655 -6343
rect 1632 -8995 1646 -6346
rect 1667 -8130 1693 -8127
rect 1667 -8159 1693 -8156
rect 1673 -8995 1687 -8159
rect 2727 -9007 2741 -3613
rect 3142 -4130 3159 -2942
rect 6646 -2944 6672 -2941
rect 4308 -2984 4340 -2981
rect 4308 -3010 4311 -2984
rect 4337 -3010 4340 -2984
rect 4308 -3013 4340 -3010
rect 5496 -3002 5522 -2999
rect 3534 -3070 3564 -3065
rect 3534 -3105 3564 -3100
rect 3542 -3131 3556 -3105
rect 3903 -3584 3929 -3581
rect 3903 -3613 3929 -3610
rect 3135 -4133 3167 -4130
rect 3135 -4159 3138 -4133
rect 3164 -4159 3167 -4133
rect 3135 -4162 3167 -4159
rect 2761 -5397 2787 -5394
rect 2761 -5426 2787 -5423
rect 2767 -9007 2781 -5426
rect 2800 -6317 2832 -6314
rect 2800 -6343 2803 -6317
rect 2829 -6343 2832 -6317
rect 2800 -6346 2832 -6343
rect 2809 -9007 2823 -6346
rect 2844 -8130 2870 -8127
rect 2844 -8159 2870 -8156
rect 2850 -9007 2864 -8159
rect 3909 -9018 3923 -3613
rect 4316 -4130 4333 -3013
rect 5496 -3031 5522 -3028
rect 4716 -3067 4746 -3062
rect 4716 -3102 4746 -3097
rect 4724 -3132 4738 -3102
rect 5089 -3584 5115 -3581
rect 5089 -3613 5115 -3610
rect 4309 -4133 4341 -4130
rect 4309 -4159 4312 -4133
rect 4338 -4159 4341 -4133
rect 4309 -4162 4341 -4159
rect 3943 -5397 3969 -5394
rect 3943 -5426 3969 -5423
rect 3949 -9018 3963 -5426
rect 3982 -6317 4014 -6314
rect 3982 -6343 3985 -6317
rect 4011 -6343 4014 -6317
rect 3982 -6346 4014 -6343
rect 3991 -9018 4005 -6346
rect 4026 -8130 4052 -8127
rect 4026 -8159 4052 -8156
rect 4032 -9018 4046 -8159
rect 5095 -9026 5109 -3613
rect 5501 -4130 5518 -3031
rect 5898 -3070 5928 -3065
rect 5898 -3105 5928 -3100
rect 5906 -3131 5920 -3105
rect 6268 -3584 6294 -3581
rect 6268 -3613 6294 -3610
rect 5497 -4133 5523 -4130
rect 5497 -4162 5523 -4159
rect 5129 -5397 5155 -5394
rect 5129 -5426 5155 -5423
rect 5135 -9026 5149 -5426
rect 5168 -6317 5200 -6314
rect 5168 -6343 5171 -6317
rect 5197 -6343 5200 -6317
rect 5168 -6346 5200 -6343
rect 5177 -9026 5191 -6346
rect 5212 -8130 5238 -8127
rect 5212 -8159 5238 -8156
rect 5218 -9026 5232 -8159
rect 6274 -9023 6288 -3613
rect 6651 -4132 6668 -2944
rect 7080 -3070 7110 -3065
rect 7080 -3105 7110 -3100
rect 7088 -3131 7102 -3105
rect 7456 -3584 7482 -3581
rect 7456 -3613 7482 -3610
rect 6647 -4135 6673 -4132
rect 6647 -4164 6673 -4161
rect 6308 -5397 6334 -5394
rect 6308 -5426 6334 -5423
rect 6314 -9023 6328 -5426
rect 6347 -6317 6379 -6314
rect 6347 -6343 6350 -6317
rect 6376 -6343 6379 -6317
rect 6347 -6346 6379 -6343
rect 6356 -9023 6370 -6346
rect 6391 -8130 6417 -8127
rect 6391 -8159 6417 -8156
rect 6397 -9023 6411 -8159
rect 7462 -9012 7476 -3613
rect 7853 -4132 7870 -2864
rect 8262 -3068 8292 -3063
rect 8262 -3103 8292 -3098
rect 8270 -3131 8284 -3103
rect 8629 -3584 8655 -3581
rect 8629 -3613 8655 -3610
rect 7849 -4135 7875 -4132
rect 7849 -4164 7875 -4161
rect 7496 -5397 7522 -5394
rect 7496 -5426 7522 -5423
rect 7502 -9012 7516 -5426
rect 7535 -6317 7567 -6314
rect 7535 -6343 7538 -6317
rect 7564 -6343 7567 -6317
rect 7535 -6346 7567 -6343
rect 7544 -9012 7558 -6346
rect 7579 -8130 7605 -8127
rect 7579 -8159 7605 -8156
rect 7585 -9012 7599 -8159
rect 8635 -9027 8649 -3613
rect 9041 -4135 9058 -2789
rect 9446 -3069 9476 -3064
rect 9446 -3104 9476 -3099
rect 9454 -3132 9468 -3104
rect 9811 -3584 9837 -3581
rect 9811 -3613 9837 -3610
rect 9034 -4161 9037 -4135
rect 9063 -4161 9066 -4135
rect 8669 -5397 8695 -5394
rect 8669 -5426 8695 -5423
rect 8675 -9027 8689 -5426
rect 8708 -6317 8740 -6314
rect 8708 -6343 8711 -6317
rect 8737 -6343 8740 -6317
rect 8708 -6346 8740 -6343
rect 8717 -9027 8731 -6346
rect 8752 -8130 8778 -8127
rect 8752 -8159 8778 -8156
rect 8758 -9027 8772 -8159
rect 9817 -9035 9831 -3613
rect 10215 -4132 10232 -2726
rect 10630 -3070 10660 -3065
rect 10630 -3105 10660 -3100
rect 10638 -3133 10652 -3105
rect 11000 -3584 11026 -3581
rect 11000 -3613 11026 -3610
rect 10211 -4135 10237 -4132
rect 10211 -4164 10237 -4161
rect 9851 -5397 9877 -5394
rect 9851 -5426 9877 -5423
rect 9857 -9035 9871 -5426
rect 9890 -6317 9922 -6314
rect 9890 -6343 9893 -6317
rect 9919 -6343 9922 -6317
rect 9890 -6346 9922 -6343
rect 9899 -9035 9913 -6346
rect 9934 -8130 9960 -8127
rect 9934 -8159 9960 -8156
rect 9940 -9035 9954 -8159
rect 11006 -9017 11020 -3613
rect 11428 -4131 11445 -2663
rect 11817 -3066 11847 -3061
rect 11817 -3101 11847 -3096
rect 11825 -3131 11839 -3101
rect 12195 -3584 12221 -3581
rect 12195 -3613 12221 -3610
rect 11424 -4134 11450 -4131
rect 11424 -4163 11450 -4160
rect 11040 -5397 11066 -5394
rect 11040 -5426 11066 -5423
rect 11046 -9017 11060 -5426
rect 11079 -6317 11111 -6314
rect 11079 -6343 11082 -6317
rect 11108 -6343 11111 -6317
rect 11079 -6346 11111 -6343
rect 11088 -9017 11102 -6346
rect 11123 -8130 11149 -8127
rect 11123 -8159 11149 -8156
rect 11129 -9017 11143 -8159
rect 12201 -9013 12215 -3613
rect 12591 -4132 12608 -2613
rect 13004 -3068 13034 -3063
rect 13004 -3103 13034 -3098
rect 13012 -3132 13026 -3103
rect 13371 -3584 13397 -3581
rect 13371 -3613 13397 -3610
rect 12587 -4135 12613 -4132
rect 12587 -4164 12613 -4161
rect 12235 -5397 12261 -5394
rect 12235 -5426 12261 -5423
rect 12241 -9013 12255 -5426
rect 12274 -6317 12306 -6314
rect 12274 -6343 12277 -6317
rect 12303 -6343 12306 -6317
rect 12274 -6346 12306 -6343
rect 12283 -9013 12297 -6346
rect 12318 -8130 12344 -8127
rect 12318 -8159 12344 -8156
rect 12324 -9013 12338 -8159
rect 13377 -9007 13391 -3613
rect 13537 -4134 13554 -2566
rect 13905 -3070 13935 -3065
rect 13905 -3105 13935 -3100
rect 13913 -3131 13927 -3105
rect 14275 -3584 14301 -3581
rect 14275 -3613 14301 -3610
rect 13530 -4160 13533 -4134
rect 13559 -4160 13562 -4134
rect 13411 -5397 13437 -5394
rect 13411 -5426 13437 -5423
rect 13417 -9007 13431 -5426
rect 13450 -6317 13482 -6314
rect 13450 -6343 13453 -6317
rect 13479 -6343 13482 -6317
rect 13450 -6346 13482 -6343
rect 13459 -9007 13473 -6346
rect 13494 -8130 13520 -8127
rect 13494 -8159 13520 -8156
rect 13500 -9007 13514 -8159
rect 14281 -9011 14295 -3613
rect 14446 -4445 14472 -4442
rect 14446 -4474 14472 -4471
rect 14315 -5397 14341 -5394
rect 14315 -5426 14341 -5423
rect 14321 -9011 14335 -5426
rect 14354 -6317 14386 -6314
rect 14354 -6343 14357 -6317
rect 14383 -6343 14386 -6317
rect 14354 -6346 14386 -6343
rect 14363 -9011 14377 -6346
rect 14398 -8130 14424 -8127
rect 14398 -8159 14424 -8156
rect 14404 -9011 14418 -8159
rect 14451 -9010 14468 -4474
rect 14502 -4534 14528 -4531
rect 14502 -4563 14528 -4560
rect 14507 -9010 14524 -4563
rect 14556 -7171 14582 -7168
rect 14556 -7200 14582 -7197
rect 14561 -9010 14578 -7200
rect 14611 -7268 14637 -7265
rect 14611 -7297 14637 -7294
rect 14616 -9010 14633 -7297
<< via2 >>
rect -4314 5031 -4284 5061
rect -4180 -2064 -4150 -2034
rect -35 -2032 -5 -2030
rect -35 -2058 -33 -2032
rect -33 -2058 -7 -2032
rect -7 -2058 -5 -2032
rect -35 -2060 -5 -2058
rect -4314 -3093 -4284 -3063
rect 524 5039 554 5069
rect 596 -637 626 -607
rect 1100 5039 1130 5069
rect 1171 -764 1201 -734
rect 1675 5039 1705 5069
rect 1751 -901 1781 -871
rect 2248 5039 2278 5069
rect 2321 -1018 2351 -988
rect 2824 5039 2854 5069
rect 2896 -1143 2926 -1113
rect 3398 5039 3428 5069
rect 3471 -1288 3501 -1258
rect 3973 5039 4003 5069
rect 4045 -1382 4075 -1380
rect 4045 -1408 4047 -1382
rect 4047 -1408 4073 -1382
rect 4073 -1408 4075 -1382
rect 4045 -1410 4075 -1408
rect 4548 5039 4578 5069
rect 4621 -1498 4651 -1468
rect 5123 5039 5153 5069
rect 5196 -1581 5226 -1551
rect 5699 5039 5729 5069
rect 5771 -1659 5801 -1629
rect 6274 5038 6304 5068
rect 6346 -1745 6376 -1715
rect 6848 5039 6878 5069
rect 6921 -1825 6951 -1795
rect 7423 5039 7453 5069
rect 7496 -1905 7526 -1875
rect 7998 5039 8028 5069
rect 8071 -1970 8101 -1940
rect 8572 5039 8602 5069
rect 8646 -2084 8676 -2054
rect 9147 5039 9177 5069
rect 9221 -2173 9251 -2143
rect 811 -2322 841 -2320
rect 811 -2348 813 -2322
rect 813 -2348 839 -2322
rect 839 -2348 841 -2322
rect 811 -2350 841 -2348
rect 1960 -2323 1990 -2321
rect 1960 -2349 1962 -2323
rect 1962 -2349 1988 -2323
rect 1988 -2349 1990 -2323
rect 1960 -2351 1990 -2349
rect 3103 -2324 3133 -2322
rect 3103 -2350 3105 -2324
rect 3105 -2350 3131 -2324
rect 3131 -2350 3133 -2324
rect 3103 -2352 3133 -2350
rect 4260 -2325 4290 -2323
rect 4260 -2351 4262 -2325
rect 4262 -2351 4288 -2325
rect 4288 -2351 4290 -2325
rect 4260 -2353 4290 -2351
rect 5400 -2323 5430 -2321
rect 5400 -2349 5402 -2323
rect 5402 -2349 5428 -2323
rect 5428 -2349 5430 -2323
rect 5400 -2351 5430 -2349
rect 6568 -2323 6598 -2321
rect 6568 -2349 6570 -2323
rect 6570 -2349 6596 -2323
rect 6596 -2349 6598 -2323
rect 6568 -2351 6598 -2349
rect 7713 -2323 7743 -2321
rect 7713 -2349 7715 -2323
rect 7715 -2349 7741 -2323
rect 7741 -2349 7743 -2323
rect 7713 -2351 7743 -2349
rect 8870 -2321 8900 -2319
rect 8870 -2347 8872 -2321
rect 8872 -2347 8898 -2321
rect 8898 -2347 8900 -2321
rect 8870 -2349 8900 -2347
rect 735 -2421 765 -2419
rect 735 -2447 737 -2421
rect 737 -2447 763 -2421
rect 763 -2447 765 -2421
rect 735 -2449 765 -2447
rect 890 -2421 920 -2419
rect 890 -2447 892 -2421
rect 892 -2447 918 -2421
rect 918 -2447 920 -2421
rect 890 -2449 920 -2447
rect 1885 -2421 1915 -2419
rect 1885 -2447 1887 -2421
rect 1887 -2447 1913 -2421
rect 1913 -2447 1915 -2421
rect 1885 -2449 1915 -2447
rect 2040 -2421 2070 -2419
rect 2040 -2447 2042 -2421
rect 2042 -2447 2068 -2421
rect 2068 -2447 2070 -2421
rect 2040 -2449 2070 -2447
rect 3035 -2421 3065 -2419
rect 3035 -2447 3037 -2421
rect 3037 -2447 3063 -2421
rect 3063 -2447 3065 -2421
rect 3035 -2449 3065 -2447
rect 3189 -2421 3219 -2419
rect 3189 -2447 3191 -2421
rect 3191 -2447 3217 -2421
rect 3217 -2447 3219 -2421
rect 3189 -2449 3219 -2447
rect 4182 -2421 4212 -2419
rect 4182 -2447 4184 -2421
rect 4184 -2447 4210 -2421
rect 4210 -2447 4212 -2421
rect 4182 -2449 4212 -2447
rect 4341 -2422 4371 -2420
rect 4341 -2448 4343 -2422
rect 4343 -2448 4369 -2422
rect 4369 -2448 4371 -2422
rect 4341 -2450 4371 -2448
rect 5334 -2421 5364 -2419
rect 5334 -2447 5336 -2421
rect 5336 -2447 5362 -2421
rect 5362 -2447 5364 -2421
rect 5334 -2449 5364 -2447
rect 5489 -2421 5519 -2419
rect 5489 -2447 5491 -2421
rect 5491 -2447 5517 -2421
rect 5517 -2447 5519 -2421
rect 5489 -2449 5519 -2447
rect 6485 -2422 6515 -2420
rect 6485 -2448 6487 -2422
rect 6487 -2448 6513 -2422
rect 6513 -2448 6515 -2422
rect 6485 -2450 6515 -2448
rect 6638 -2422 6668 -2420
rect 6638 -2448 6640 -2422
rect 6640 -2448 6666 -2422
rect 6666 -2448 6668 -2422
rect 6638 -2450 6668 -2448
rect 7636 -2421 7666 -2419
rect 7636 -2447 7638 -2421
rect 7638 -2447 7664 -2421
rect 7664 -2447 7666 -2421
rect 7636 -2449 7666 -2447
rect 7789 -2421 7819 -2419
rect 7789 -2447 7791 -2421
rect 7791 -2447 7817 -2421
rect 7817 -2447 7819 -2421
rect 7789 -2449 7819 -2447
rect 8785 -2420 8815 -2418
rect 8785 -2446 8787 -2420
rect 8787 -2446 8813 -2420
rect 8813 -2446 8815 -2420
rect 8785 -2448 8815 -2446
rect 8937 -2421 8967 -2419
rect 8937 -2447 8939 -2421
rect 8939 -2447 8965 -2421
rect 8965 -2447 8967 -2421
rect 8937 -2449 8967 -2447
rect 466 -2498 496 -2496
rect 466 -2524 468 -2498
rect 468 -2524 494 -2498
rect 494 -2524 496 -2498
rect 466 -2526 496 -2524
rect 1159 -2491 1189 -2489
rect 1159 -2517 1161 -2491
rect 1161 -2517 1187 -2491
rect 1187 -2517 1189 -2491
rect 1159 -2519 1189 -2517
rect 1615 -2490 1645 -2488
rect 1615 -2516 1617 -2490
rect 1617 -2516 1643 -2490
rect 1643 -2516 1645 -2490
rect 1615 -2518 1645 -2516
rect 2308 -2495 2338 -2493
rect 2308 -2521 2310 -2495
rect 2310 -2521 2336 -2495
rect 2336 -2521 2338 -2495
rect 2308 -2523 2338 -2521
rect 2767 -2496 2797 -2494
rect 2767 -2522 2769 -2496
rect 2769 -2522 2795 -2496
rect 2795 -2522 2797 -2496
rect 2767 -2524 2797 -2522
rect 3459 -2494 3489 -2492
rect 3459 -2520 3461 -2494
rect 3461 -2520 3487 -2494
rect 3487 -2520 3489 -2494
rect 3459 -2522 3489 -2520
rect 3917 -2496 3947 -2494
rect 3917 -2522 3919 -2496
rect 3919 -2522 3945 -2496
rect 3945 -2522 3947 -2496
rect 3917 -2524 3947 -2522
rect 4608 -2498 4638 -2496
rect 4608 -2524 4610 -2498
rect 4610 -2524 4636 -2498
rect 4636 -2524 4638 -2498
rect 4608 -2526 4638 -2524
rect 5066 -2492 5096 -2490
rect 5066 -2518 5068 -2492
rect 5068 -2518 5094 -2492
rect 5094 -2518 5096 -2492
rect 5066 -2520 5096 -2518
rect 5759 -2494 5789 -2492
rect 5759 -2520 5761 -2494
rect 5761 -2520 5787 -2494
rect 5787 -2520 5789 -2494
rect 5759 -2522 5789 -2520
rect 6216 -2490 6246 -2488
rect 6216 -2516 6218 -2490
rect 6218 -2516 6244 -2490
rect 6244 -2516 6246 -2490
rect 6216 -2518 6246 -2516
rect 6908 -2494 6938 -2492
rect 6908 -2520 6910 -2494
rect 6910 -2520 6936 -2494
rect 6936 -2520 6938 -2494
rect 6908 -2522 6938 -2520
rect 7366 -2494 7396 -2492
rect 7366 -2520 7368 -2494
rect 7368 -2520 7394 -2494
rect 7394 -2520 7396 -2494
rect 7366 -2522 7396 -2520
rect 8058 -2497 8088 -2495
rect 8058 -2523 8060 -2497
rect 8060 -2523 8086 -2497
rect 8086 -2523 8088 -2497
rect 8058 -2525 8088 -2523
rect 8516 -2495 8546 -2493
rect 8516 -2521 8518 -2495
rect 8518 -2521 8544 -2495
rect 8544 -2521 8546 -2495
rect 8516 -2523 8546 -2521
rect 9207 -2520 9235 -2492
rect -3524 -3097 -3494 -3067
rect -2374 -3097 -2344 -3067
rect -1192 -3096 -1162 -3066
rect -11 -3101 19 -3071
rect 1170 -3099 1200 -3069
rect 2352 -3100 2382 -3070
rect 3534 -3100 3564 -3070
rect 4716 -3097 4746 -3067
rect 5898 -3100 5928 -3070
rect 7080 -3100 7110 -3070
rect 8262 -3098 8292 -3068
rect 9446 -3099 9476 -3069
rect 10630 -3100 10660 -3070
rect 11817 -3096 11847 -3066
rect 13004 -3098 13034 -3068
rect 13905 -3100 13935 -3070
<< metal3 >>
rect 519 5069 559 5074
rect 519 5064 524 5069
rect -4549 5061 524 5064
rect -4549 5034 -4314 5061
rect -4317 5031 -4314 5034
rect -4284 5039 524 5061
rect 554 5064 559 5069
rect 1095 5069 1135 5074
rect 1095 5064 1100 5069
rect 554 5039 1100 5064
rect 1130 5064 1135 5069
rect 1670 5069 1710 5074
rect 1670 5064 1675 5069
rect 1130 5039 1675 5064
rect 1705 5064 1710 5069
rect 2243 5069 2283 5074
rect 2243 5064 2248 5069
rect 1705 5039 2248 5064
rect 2278 5064 2283 5069
rect 2819 5069 2859 5074
rect 2819 5064 2824 5069
rect 2278 5039 2824 5064
rect 2854 5064 2859 5069
rect 3393 5069 3433 5074
rect 3393 5064 3398 5069
rect 2854 5039 3398 5064
rect 3428 5064 3433 5069
rect 3968 5069 4008 5074
rect 3968 5064 3973 5069
rect 3428 5039 3973 5064
rect 4003 5064 4008 5069
rect 4543 5069 4583 5074
rect 4543 5064 4548 5069
rect 4003 5039 4548 5064
rect 4578 5064 4583 5069
rect 5118 5069 5158 5074
rect 5118 5064 5123 5069
rect 4578 5039 5123 5064
rect 5153 5064 5158 5069
rect 5694 5069 5734 5074
rect 5694 5064 5699 5069
rect 5153 5039 5699 5064
rect 5729 5064 5734 5069
rect 6269 5068 6309 5073
rect 6269 5064 6274 5068
rect 5729 5039 6274 5064
rect -4284 5038 6274 5039
rect 6304 5064 6309 5068
rect 6843 5069 6883 5074
rect 6843 5064 6848 5069
rect 6304 5039 6848 5064
rect 6878 5064 6883 5069
rect 7418 5069 7458 5074
rect 7418 5064 7423 5069
rect 6878 5039 7423 5064
rect 7453 5064 7458 5069
rect 7993 5069 8033 5074
rect 7993 5064 7998 5069
rect 7453 5039 7998 5064
rect 8028 5064 8033 5069
rect 8567 5069 8607 5074
rect 8567 5064 8572 5069
rect 8028 5039 8572 5064
rect 8602 5064 8607 5069
rect 9142 5069 9182 5074
rect 9142 5064 9147 5069
rect 8602 5039 9147 5064
rect 9177 5064 9182 5069
rect 9177 5039 10038 5064
rect 6304 5038 10038 5039
rect -4284 5034 10038 5038
rect -4284 5031 -4281 5034
rect 6269 5033 6309 5034
rect -4317 5028 -4281 5031
rect 593 -607 629 -604
rect 593 -637 596 -607
rect 626 -637 10048 -607
rect 593 -640 629 -637
rect 1168 -734 1204 -731
rect 1168 -764 1171 -734
rect 1201 -764 10048 -734
rect 1168 -767 1204 -764
rect 1748 -871 1784 -868
rect 1748 -901 1751 -871
rect 1781 -901 10048 -871
rect 1748 -904 1784 -901
rect 2318 -988 2354 -985
rect 2318 -1018 2321 -988
rect 2351 -1018 10048 -988
rect 2318 -1021 2354 -1018
rect 2893 -1113 2929 -1110
rect 2893 -1143 2896 -1113
rect 2926 -1143 10048 -1113
rect 2893 -1146 2929 -1143
rect 3468 -1258 3504 -1255
rect 3468 -1288 3471 -1258
rect 3501 -1288 10048 -1258
rect 3468 -1291 3504 -1288
rect 4040 -1380 4080 -1375
rect 4040 -1410 4045 -1380
rect 4075 -1410 10048 -1380
rect 4040 -1415 4080 -1410
rect 4618 -1468 4654 -1465
rect 4618 -1498 4621 -1468
rect 4651 -1498 10048 -1468
rect 4618 -1501 4654 -1498
rect 5193 -1551 5229 -1548
rect 5193 -1581 5196 -1551
rect 5226 -1581 10048 -1551
rect 5193 -1584 5229 -1581
rect 5768 -1629 5804 -1626
rect 5768 -1659 5771 -1629
rect 5801 -1659 10048 -1629
rect 5768 -1662 5804 -1659
rect 6343 -1715 6379 -1712
rect 6343 -1745 6346 -1715
rect 6376 -1745 10048 -1715
rect 6343 -1748 6379 -1745
rect 6918 -1795 6954 -1792
rect 6918 -1825 6921 -1795
rect 6951 -1825 10048 -1795
rect 6918 -1828 6954 -1825
rect 7493 -1875 7529 -1872
rect 7493 -1905 7496 -1875
rect 7526 -1905 10048 -1875
rect 7493 -1908 7529 -1905
rect 8068 -1940 8104 -1937
rect 8068 -1970 8071 -1940
rect 8101 -1970 10048 -1940
rect 8068 -1973 8104 -1970
rect -40 -2030 0 -2025
rect -4552 -2034 -35 -2030
rect -4552 -2060 -4180 -2034
rect -4183 -2064 -4180 -2060
rect -4150 -2060 -35 -2034
rect -5 -2060 0 -2030
rect -4150 -2064 -4147 -2060
rect -4183 -2067 -4147 -2064
rect -40 -2065 0 -2060
rect 8643 -2054 8679 -2051
rect -35 -2321 -5 -2065
rect 8643 -2084 8646 -2054
rect 8676 -2084 10048 -2054
rect 8643 -2087 8679 -2084
rect 9218 -2143 9254 -2140
rect 9218 -2173 9221 -2143
rect 9251 -2173 10048 -2143
rect 9218 -2176 9254 -2173
rect 806 -2320 846 -2315
rect 805 -2321 811 -2320
rect -35 -2350 811 -2321
rect 841 -2321 846 -2320
rect 1955 -2321 1995 -2316
rect 3098 -2321 3138 -2317
rect 4255 -2321 4295 -2318
rect 5395 -2321 5435 -2316
rect 6563 -2321 6603 -2316
rect 7708 -2321 7748 -2316
rect 8865 -2319 8905 -2314
rect 8864 -2321 8870 -2319
rect 841 -2350 1960 -2321
rect -35 -2351 1960 -2350
rect 1990 -2322 5400 -2321
rect 1990 -2351 3103 -2322
rect 806 -2355 846 -2351
rect 1955 -2356 1995 -2351
rect 3097 -2352 3103 -2351
rect 3133 -2323 5400 -2322
rect 3133 -2351 4260 -2323
rect 3133 -2352 3138 -2351
rect 3098 -2357 3138 -2352
rect 4254 -2353 4260 -2351
rect 4290 -2351 5400 -2323
rect 5430 -2351 6568 -2321
rect 6598 -2351 7713 -2321
rect 7743 -2349 8870 -2321
rect 8900 -2349 8905 -2319
rect 7743 -2351 8905 -2349
rect 4290 -2353 4295 -2351
rect 4255 -2358 4295 -2353
rect 5395 -2356 5435 -2351
rect 6563 -2356 6603 -2351
rect 7708 -2356 7748 -2351
rect 8865 -2354 8905 -2351
rect 730 -2419 770 -2414
rect 885 -2419 925 -2414
rect 1880 -2419 1920 -2414
rect 2035 -2419 2075 -2414
rect 3030 -2419 3070 -2414
rect 3184 -2419 3224 -2414
rect 4177 -2419 4217 -2414
rect 4336 -2419 4376 -2415
rect 5329 -2419 5369 -2414
rect 5484 -2419 5524 -2414
rect 6480 -2419 6520 -2415
rect 6633 -2419 6673 -2415
rect 7631 -2419 7671 -2414
rect 7784 -2419 7824 -2414
rect 8780 -2418 8820 -2414
rect 8780 -2419 8785 -2418
rect -4542 -2449 735 -2419
rect 765 -2449 890 -2419
rect 920 -2449 1885 -2419
rect 1915 -2449 2040 -2419
rect 2070 -2449 3035 -2419
rect 3065 -2449 3189 -2419
rect 3219 -2449 4182 -2419
rect 4212 -2420 5334 -2419
rect 4212 -2449 4341 -2420
rect 730 -2454 770 -2449
rect 885 -2454 925 -2449
rect 1880 -2454 1920 -2449
rect 2035 -2454 2075 -2449
rect 3030 -2454 3070 -2449
rect 3184 -2454 3224 -2449
rect 4177 -2454 4217 -2449
rect 4336 -2450 4341 -2449
rect 4371 -2449 5334 -2420
rect 5364 -2449 5489 -2419
rect 5519 -2420 7636 -2419
rect 5519 -2449 6485 -2420
rect 4371 -2450 4376 -2449
rect 4336 -2455 4376 -2450
rect 5329 -2454 5369 -2449
rect 5484 -2454 5524 -2449
rect 6480 -2450 6485 -2449
rect 6515 -2449 6638 -2420
rect 6515 -2450 6520 -2449
rect 6480 -2455 6520 -2450
rect 6633 -2450 6638 -2449
rect 6668 -2449 7636 -2420
rect 7666 -2449 7789 -2419
rect 7819 -2448 8785 -2419
rect 8815 -2419 8820 -2418
rect 8932 -2419 8972 -2413
rect 8815 -2448 8937 -2419
rect 7819 -2449 8937 -2448
rect 8967 -2449 8972 -2419
rect 6668 -2450 6673 -2449
rect 6633 -2455 6673 -2450
rect 7631 -2454 7671 -2449
rect 7784 -2454 7824 -2449
rect 8780 -2454 8820 -2449
rect 8932 -2454 8972 -2449
rect 1154 -2489 1194 -2484
rect 461 -2495 501 -2491
rect 1154 -2495 1159 -2489
rect -4542 -2496 1159 -2495
rect -4542 -2525 466 -2496
rect 461 -2526 466 -2525
rect 496 -2519 1159 -2496
rect 1189 -2495 1194 -2489
rect 1610 -2488 1650 -2483
rect 1610 -2495 1615 -2488
rect 1189 -2518 1615 -2495
rect 1645 -2495 1650 -2488
rect 2303 -2493 2343 -2488
rect 2303 -2495 2308 -2493
rect 1645 -2518 2308 -2495
rect 1189 -2519 2308 -2518
rect 496 -2523 2308 -2519
rect 2338 -2495 2343 -2493
rect 2762 -2494 2802 -2489
rect 2762 -2495 2767 -2494
rect 2338 -2523 2767 -2495
rect 496 -2524 2767 -2523
rect 2797 -2495 2802 -2494
rect 3454 -2492 3494 -2487
rect 3454 -2495 3459 -2492
rect 2797 -2522 3459 -2495
rect 3489 -2495 3494 -2492
rect 3912 -2494 3952 -2489
rect 5061 -2490 5101 -2485
rect 3912 -2495 3917 -2494
rect 3489 -2522 3917 -2495
rect 2797 -2524 3917 -2522
rect 3947 -2495 3952 -2494
rect 4603 -2495 4643 -2491
rect 5061 -2495 5066 -2490
rect 3947 -2496 5066 -2495
rect 3947 -2524 4608 -2496
rect 496 -2525 4608 -2524
rect 496 -2526 501 -2525
rect 461 -2531 501 -2526
rect 2303 -2528 2343 -2525
rect 2762 -2529 2802 -2525
rect 3454 -2527 3494 -2525
rect 3912 -2529 3952 -2525
rect 4603 -2526 4608 -2525
rect 4638 -2520 5066 -2496
rect 5096 -2495 5101 -2490
rect 5754 -2492 5794 -2487
rect 5754 -2495 5759 -2492
rect 5096 -2520 5759 -2495
rect 4638 -2522 5759 -2520
rect 5789 -2495 5794 -2492
rect 6211 -2488 6251 -2483
rect 6211 -2495 6216 -2488
rect 5789 -2518 6216 -2495
rect 6246 -2495 6251 -2488
rect 6903 -2492 6943 -2487
rect 6903 -2495 6908 -2492
rect 6246 -2518 6908 -2495
rect 5789 -2522 6908 -2518
rect 6938 -2495 6943 -2492
rect 7361 -2492 7401 -2487
rect 7361 -2495 7366 -2492
rect 6938 -2522 7366 -2495
rect 7396 -2495 7401 -2492
rect 8053 -2495 8093 -2490
rect 8511 -2493 8551 -2489
rect 8511 -2495 8516 -2493
rect 7396 -2522 8058 -2495
rect 4638 -2525 8058 -2522
rect 8088 -2523 8516 -2495
rect 8546 -2495 8551 -2493
rect 9203 -2492 9239 -2487
rect 9203 -2495 9207 -2492
rect 8546 -2520 9207 -2495
rect 9235 -2520 9239 -2492
rect 8546 -2523 9239 -2520
rect 8088 -2525 9239 -2523
rect 4638 -2526 4643 -2525
rect 4603 -2531 4643 -2526
rect 5754 -2527 5794 -2525
rect 6903 -2527 6943 -2525
rect 7361 -2527 7401 -2525
rect 8053 -2530 8093 -2525
rect 8511 -2529 8551 -2525
rect -4317 -3063 -4281 -3060
rect -4317 -3067 -4314 -3063
rect -4515 -3093 -4314 -3067
rect -4284 -3067 -4281 -3063
rect -3527 -3067 -3491 -3064
rect -2377 -3067 -2341 -3064
rect -1195 -3066 -1159 -3063
rect -1195 -3067 -1192 -3066
rect -4284 -3093 -3524 -3067
rect -4515 -3097 -3524 -3093
rect -3494 -3097 -2374 -3067
rect -2344 -3096 -1192 -3067
rect -1162 -3067 -1159 -3066
rect 1167 -3067 1203 -3066
rect 4713 -3067 4749 -3064
rect 8259 -3067 8295 -3065
rect 11814 -3066 11850 -3063
rect 9443 -3067 9479 -3066
rect 11814 -3067 11817 -3066
rect -1162 -3069 4716 -3067
rect -1162 -3071 1170 -3069
rect -1162 -3096 -11 -3071
rect -2344 -3097 -11 -3096
rect -3527 -3100 -3491 -3097
rect -2377 -3100 -2341 -3097
rect -1195 -3099 -1159 -3097
rect -14 -3101 -11 -3097
rect 19 -3097 1170 -3071
rect 19 -3101 22 -3097
rect -14 -3104 22 -3101
rect 1167 -3099 1170 -3097
rect 1200 -3070 4716 -3069
rect 1200 -3097 2352 -3070
rect 1200 -3099 1203 -3097
rect 1167 -3102 1203 -3099
rect 2349 -3100 2352 -3097
rect 2382 -3097 3534 -3070
rect 2382 -3100 2385 -3097
rect 2349 -3103 2385 -3100
rect 3531 -3100 3534 -3097
rect 3564 -3097 4716 -3070
rect 4746 -3068 11817 -3067
rect 4746 -3070 8262 -3068
rect 4746 -3097 5898 -3070
rect 3564 -3100 3567 -3097
rect 4713 -3100 4749 -3097
rect 5895 -3100 5898 -3097
rect 5928 -3097 7080 -3070
rect 5928 -3100 5931 -3097
rect 3531 -3103 3567 -3100
rect 5895 -3103 5931 -3100
rect 7077 -3100 7080 -3097
rect 7110 -3097 8262 -3070
rect 7110 -3100 7113 -3097
rect 7077 -3103 7113 -3100
rect 8259 -3098 8262 -3097
rect 8292 -3069 11817 -3068
rect 8292 -3097 9446 -3069
rect 8292 -3098 8295 -3097
rect 8259 -3101 8295 -3098
rect 9443 -3099 9446 -3097
rect 9476 -3070 11817 -3069
rect 9476 -3097 10630 -3070
rect 9476 -3099 9479 -3097
rect 9443 -3102 9479 -3099
rect 10627 -3100 10630 -3097
rect 10660 -3096 11817 -3070
rect 11847 -3067 11850 -3066
rect 13001 -3067 13037 -3065
rect 11847 -3068 14436 -3067
rect 11847 -3096 13004 -3068
rect 10660 -3097 13004 -3096
rect 10660 -3100 10663 -3097
rect 11814 -3099 11850 -3097
rect 13001 -3098 13004 -3097
rect 13034 -3070 14436 -3068
rect 13034 -3097 13905 -3070
rect 13034 -3098 13037 -3097
rect 10627 -3103 10663 -3100
rect 13001 -3101 13037 -3098
rect 13902 -3100 13905 -3097
rect 13935 -3097 14436 -3070
rect 13935 -3100 13938 -3097
rect 13902 -3103 13938 -3100
use 1  1_0
timestamp 1661016133
transform 1 0 225 0 1 3818
box 0 0 9241 270
use 1  1_1
timestamp 1661016133
transform 1 0 225 0 1 4356
box 0 0 9241 270
use 1  1_2
timestamp 1661016133
transform 1 0 225 0 1 4597
box 0 0 9241 270
use 1  1_3
timestamp 1661016133
transform 1 0 225 0 1 -360
box 0 0 9241 270
use 1  1_4
timestamp 1661016133
transform 1 0 225 0 1 -601
box 0 0 9241 270
use 1  1_5
timestamp 1661016133
transform 1 0 225 0 1 -1142
box 0 0 9241 270
use 3  3_0
timestamp 1661016133
transform 1 0 1047 0 1 3849
box -822 210 8419 480
use 3  3_1
timestamp 1661016133
transform 1 0 1047 0 1 -1111
box -822 210 8419 480
use ADC_vertical  ADC_vertical_0
timestamp 1662726195
transform 1 0 -3212 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_1
timestamp 1662726195
transform 1 0 -2031 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_2
timestamp 1662726195
transform 1 0 -849 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_3
timestamp 1662726195
transform 1 0 333 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_4
timestamp 1662726195
transform 1 0 1515 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_5
timestamp 1662726195
transform 1 0 2697 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_6
timestamp 1662726195
transform 1 0 3879 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_7
timestamp 1662726195
transform 1 0 5061 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_8
timestamp 1662726195
transform 1 0 6245 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_9
timestamp 1662726195
transform 1 0 7429 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_10
timestamp 1662726195
transform 1 0 8616 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_11
timestamp 1662726195
transform 1 0 9803 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_12
timestamp 1662726195
transform 1 0 10704 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_13
timestamp 1662726195
transform 1 0 -4393 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_14
timestamp 1662726195
transform 1 0 -5575 0 1 -3254
box 2881 -5370 3543 137
use ADC_vertical  ADC_vertical_15
timestamp 1662726195
transform 1 0 -6725 0 1 -3254
box 2881 -5370 3543 137
use Array_16x16  Array_16x16_0
timestamp 1661018830
transform 1 0 -151 0 1 3625
box 376 -3744 9617 222
use Precharge  Precharge_0
timestamp 1661012742
transform 1 0 -996 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_1
timestamp 1661012742
transform 1 0 -421 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_2
timestamp 1661012742
transform 1 0 154 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_3
timestamp 1661012742
transform 1 0 729 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_4
timestamp 1661012742
transform 1 0 1304 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_5
timestamp 1661012742
transform 1 0 1879 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_6
timestamp 1661012742
transform 1 0 2454 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_7
timestamp 1661012742
transform 1 0 3029 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_8
timestamp 1661012742
transform 1 0 3604 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_9
timestamp 1661012742
transform 1 0 4179 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_10
timestamp 1661012742
transform 1 0 4754 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_11
timestamp 1661012742
transform 1 0 5329 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_12
timestamp 1661012742
transform 1 0 5904 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_13
timestamp 1661012742
transform 1 0 6479 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_14
timestamp 1661012742
transform 1 0 7054 0 1 4697
box 1221 170 1837 362
use Precharge  Precharge_15
timestamp 1661012742
transform 1 0 7629 0 1 4697
box 1221 170 1837 362
use Sense_amplifier  Sense_amplifier_0
timestamp 1662579941
transform 1 0 -1547 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_1
timestamp 1662579941
transform 1 0 -972 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_2
timestamp 1662579941
transform 1 0 -397 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_3
timestamp 1662579941
transform 1 0 178 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_4
timestamp 1662579941
transform 1 0 753 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_5
timestamp 1662579941
transform 1 0 1328 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_6
timestamp 1662579941
transform 1 0 1903 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_7
timestamp 1662579941
transform 1 0 2478 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_8
timestamp 1662579941
transform 1 0 3053 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_9
timestamp 1662579941
transform 1 0 3628 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_10
timestamp 1662579941
transform 1 0 4203 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_11
timestamp 1662579941
transform 1 0 4778 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_12
timestamp 1662579941
transform 1 0 5353 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_13
timestamp 1662579941
transform 1 0 5928 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_14
timestamp 1662579941
transform 1 0 6503 0 1 -1052
box 1772 -874 2388 -90
use Sense_amplifier  Sense_amplifier_15
timestamp 1662579941
transform 1 0 7078 0 1 -1052
box 1772 -874 2388 -90
use Write_driver  Write_driver_0
timestamp 1662369180
transform 1 0 -12 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_1
timestamp 1662369180
transform 1 0 563 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_2
timestamp 1662369180
transform 1 0 1138 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_3
timestamp 1662369180
transform 1 0 1713 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_4
timestamp 1662369180
transform 1 0 2288 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_5
timestamp 1662369180
transform 1 0 2863 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_6
timestamp 1662369180
transform 1 0 3438 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_7
timestamp 1662369180
transform 1 0 4013 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_8
timestamp 1662369180
transform 1 0 4588 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_9
timestamp 1662369180
transform 1 0 5163 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_10
timestamp 1662369180
transform 1 0 5738 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_11
timestamp 1662369180
transform 1 0 6313 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_12
timestamp 1662369180
transform 1 0 6888 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_13
timestamp 1662369180
transform 1 0 7463 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_14
timestamp 1662369180
transform 1 0 8038 0 1 -1791
box 237 -465 853 -125
use Write_driver  Write_driver_15
timestamp 1662369180
transform 1 0 8613 0 1 -1791
box 237 -465 853 -125
use substrate_contact  substrate_contact_0
timestamp 1661018752
transform 1 0 -12152 0 1 4611
box 12377 -317 21618 -203
use substrate_contact  substrate_contact_1
timestamp 1661018752
transform 1 0 -12152 0 1 -346
box 12377 -317 21618 -203
<< labels >>
flabel space -3191 225 -3177 228 0 FreeSans 80 0 0 0 RWLB[2]
port 97 nsew
flabel metal2 240 5353 240 5353 0 FreeSans 40 0 0 0 Din[0]
port 263 nsew
flabel metal2 821 5342 821 5342 0 FreeSans 40 0 0 0 Din[1]
port 264 nsew
flabel metal2 1391 5339 1391 5339 0 FreeSans 40 0 0 0 Din[2]
port 265 nsew
flabel metal2 1970 5340 1970 5340 0 FreeSans 40 0 0 0 Din[3]
port 266 nsew
flabel metal2 2543 5340 2543 5340 0 FreeSans 40 0 0 0 Din[4]
port 267 nsew
flabel metal2 3116 5338 3116 5338 0 FreeSans 40 0 0 0 Din[5]
port 268 nsew
flabel metal2 3692 5339 3692 5339 0 FreeSans 40 0 0 0 Din[6]
port 269 nsew
flabel metal2 4270 5340 4270 5340 0 FreeSans 40 0 0 0 Din[7]
port 270 nsew
flabel metal2 4844 5340 4844 5340 0 FreeSans 40 0 0 0 Din[8]
port 271 nsew
flabel metal2 5418 5338 5418 5338 0 FreeSans 40 0 0 0 Din[9]
port 272 nsew
flabel metal2 5994 5339 5994 5339 0 FreeSans 40 0 0 0 Din[10]
port 273 nsew
flabel metal2 6567 5339 6567 5339 0 FreeSans 40 0 0 0 Din[11]
port 274 nsew
flabel metal2 7142 5339 7142 5339 0 FreeSans 40 0 0 0 Din[12]
port 275 nsew
flabel metal2 7718 5340 7718 5340 0 FreeSans 40 0 0 0 Din[13]
port 276 nsew
flabel metal2 8295 5340 8295 5340 0 FreeSans 40 0 0 0 Din[14]
port 277 nsew
flabel metal2 8869 5340 8869 5340 0 FreeSans 40 0 0 0 Din[15]
port 278 nsew
flabel metal1 -4549 3741 -4546 3755 0 FreeSans 80 0 0 0 RWL[0]
port 87 nsew
flabel metal1 -4549 3701 -4546 3715 0 FreeSans 80 0 0 0 WWL[0]
port 88 nsew
flabel metal1 -4549 3660 -4546 3674 0 FreeSans 80 0 0 0 RWLB[0]
port 89 nsew
flabel metal1 -4549 3500 -4546 3514 0 FreeSans 80 0 0 0 RWL[1]
port 91 nsew
flabel metal1 -4549 3460 -4546 3474 0 FreeSans 80 0 0 0 WWL[1]
port 92 nsew
flabel metal1 -4549 3419 -4546 3433 0 FreeSans 80 0 0 0 RWLB[1]
port 93 nsew
flabel metal1 -4549 3259 -4546 3273 0 FreeSans 80 0 0 0 RWL[2]
port 95 nsew
flabel metal1 -4549 3219 -4546 3233 0 FreeSans 80 0 0 0 WWL[2]
port 96 nsew
flabel metal1 -4549 3178 -4546 3192 0 FreeSans 80 0 0 0 RWLB[2]
port 98 nsew
flabel metal1 -4549 3018 -4546 3032 0 FreeSans 80 0 0 0 RWL[3]
port 100 nsew
flabel metal1 -4549 2978 -4546 2992 0 FreeSans 80 0 0 0 WWL[3]
port 101 nsew
flabel metal1 -4549 2937 -4546 2951 0 FreeSans 80 0 0 0 RWLB[3]
port 102 nsew
flabel metal1 -4549 2737 -4546 2751 0 FreeSans 80 0 0 0 RWL[4]
port 104 nsew
flabel metal1 -4549 2697 -4546 2711 0 FreeSans 80 0 0 0 WWL[4]
port 105 nsew
flabel metal1 -4549 2656 -4546 2670 0 FreeSans 80 0 0 0 RWLB[4]
port 106 nsew
flabel metal1 -4549 2496 -4546 2510 0 FreeSans 80 0 0 0 RWL[5]
port 111 nsew
flabel metal1 -4549 2456 -4546 2470 0 FreeSans 80 0 0 0 WWL[5]
port 112 nsew
flabel metal1 -4549 2415 -4546 2429 0 FreeSans 80 0 0 0 RWLB[5]
port 113 nsew
flabel metal1 -4549 2255 -4546 2269 0 FreeSans 80 0 0 0 RWL[6]
port 115 nsew
flabel metal1 -4549 2215 -4546 2229 0 FreeSans 80 0 0 0 WWL[6]
port 116 nsew
flabel metal1 -4549 2174 -4546 2188 0 FreeSans 80 0 0 0 RWLB[6]
port 117 nsew
flabel metal1 -4549 2014 -4546 2028 0 FreeSans 80 0 0 0 RWL[7]
port 119 nsew
flabel metal1 -4549 1974 -4546 1988 0 FreeSans 80 0 0 0 WWL[7]
port 120 nsew
flabel metal1 -4549 1933 -4546 1947 0 FreeSans 80 0 0 0 RWLB[7]
port 121 nsew
flabel metal1 -4549 1773 -4546 1787 0 FreeSans 80 0 0 0 RWL[8]
port 123 nsew
flabel metal1 -4549 1733 -4546 1747 0 FreeSans 80 0 0 0 WWL[8]
port 124 nsew
flabel metal1 -4549 1692 -4546 1706 0 FreeSans 80 0 0 0 RWLB[8]
port 125 nsew
flabel metal1 -4549 1532 -4546 1546 0 FreeSans 80 0 0 0 RWL[9]
port 127 nsew
flabel metal1 -4549 1492 -4546 1506 0 FreeSans 80 0 0 0 WWL[9]
port 128 nsew
flabel metal1 -4549 1451 -4546 1465 0 FreeSans 80 0 0 0 RWLB[9]
port 129 nsew
flabel metal1 -4549 1291 -4546 1305 0 FreeSans 80 0 0 0 RWL[10]
port 131 nsew
flabel metal1 -4549 1251 -4546 1265 0 FreeSans 80 0 0 0 WWL[10]
port 132 nsew
flabel metal1 -4549 1210 -4546 1224 0 FreeSans 80 0 0 0 RWLB[10]
port 133 nsew
flabel metal1 -4549 1050 -4546 1064 0 FreeSans 80 0 0 0 RWL[11]
port 135 nsew
flabel metal1 -4549 1010 -4546 1024 0 FreeSans 80 0 0 0 WWL[11]
port 136 nsew
flabel metal1 -4549 969 -4546 983 0 FreeSans 80 0 0 0 RWLB[11]
port 137 nsew
flabel metal1 -4549 768 -4546 782 0 FreeSans 80 0 0 0 RWL[12]
port 139 nsew
flabel metal1 -4549 728 -4546 742 0 FreeSans 80 0 0 0 WWL[12]
port 140 nsew
flabel metal1 -4549 687 -4546 701 0 FreeSans 80 0 0 0 RWLB[12]
port 141 nsew
flabel metal1 -4549 527 -4546 541 0 FreeSans 80 0 0 0 RWL[13]
port 143 nsew
flabel metal1 -4549 487 -4546 501 0 FreeSans 80 0 0 0 WWL[13]
port 144 nsew
flabel metal1 -4549 446 -4546 460 0 FreeSans 80 0 0 0 RWLB[13]
port 145 nsew
flabel metal1 -4549 286 -4546 300 0 FreeSans 80 0 0 0 RWL[14]
port 147 nsew
flabel metal1 -4549 246 -4546 260 0 FreeSans 80 0 0 0 WWL[14]
port 148 nsew
flabel metal1 -4549 205 -4546 219 0 FreeSans 80 0 0 0 RWLB[14]
port 149 nsew
flabel metal1 -4549 45 -4546 59 0 FreeSans 80 0 0 0 RWL[15]
port 150 nsew
flabel metal1 -4549 5 -4546 19 0 FreeSans 80 0 0 0 WWL[15]
port 152 nsew
flabel metal1 -4549 -36 -4546 -22 0 FreeSans 80 0 0 0 RWLB[15]
port 153 nsew
flabel metal1 -4549 4721 -4546 4735 0 FreeSans 80 0 0 0 WWLD[0]
port 279 nsew
flabel metal1 -4549 4480 -4546 4494 0 FreeSans 80 0 0 0 WWLD[1]
port 280 nsew
flabel metal1 -4549 4183 -4546 4197 0 FreeSans 80 0 0 0 WWLD[2]
port 281 nsew
flabel metal1 -4549 3942 -4546 3956 0 FreeSans 80 0 0 0 WWLD[3]
port 282 nsew
flabel metal1 -4549 -236 -4546 -222 0 FreeSans 80 0 0 0 WWLD[4]
port 283 nsew
flabel metal1 -4549 -477 -4546 -463 0 FreeSans 80 0 0 0 WWLD[5]
port 284 nsew
flabel metal1 -4549 -777 -4546 -763 0 FreeSans 80 0 0 0 WWLD[6]
port 285 nsew
flabel metal1 -4549 -1018 -4546 -1004 0 FreeSans 80 0 0 0 WWLD[7]
port 286 nsew
flabel metal1 -4544 -1866 -4541 -1852 0 FreeSans 80 0 0 0 PRE_VLSA
port 155 nsew
flabel metal1 -4544 -1964 -4541 -1950 0 FreeSans 80 0 0 0 WE
port 157 nsew
flabel metal3 10042 -622 10042 -622 0 FreeSans 80 0 0 0 SA_OUT[0]
port 287 nsew
flabel metal3 10032 -751 10032 -751 0 FreeSans 80 0 0 0 SA_OUT[1]
port 288 nsew
flabel metal3 10037 -886 10037 -886 0 FreeSans 80 0 0 0 SA_OUT[2]
port 289 nsew
flabel metal3 10034 -1003 10034 -1003 0 FreeSans 80 0 0 0 SA_OUT[3]
port 290 nsew
flabel metal3 10035 -1128 10035 -1128 0 FreeSans 80 0 0 0 SA_OUT[4]
port 291 nsew
flabel metal3 10034 -1274 10034 -1274 0 FreeSans 80 0 0 0 SA_OUT[5]
port 294 nsew
flabel metal3 10033 -1395 10033 -1395 0 FreeSans 80 0 0 0 SA_OUT[6]
port 295 nsew
flabel metal3 10031 -1481 10031 -1481 0 FreeSans 80 0 0 0 SA_OUT[7]
port 296 nsew
flabel metal3 10037 -1566 10037 -1566 0 FreeSans 80 0 0 0 SA_OUT[8]
port 297 nsew
flabel metal3 10034 -1644 10034 -1644 0 FreeSans 80 0 0 0 SA_OUT[9]
port 298 nsew
flabel metal3 10030 -1731 10030 -1731 0 FreeSans 80 0 0 0 SA_OUT[10]
port 299 nsew
flabel metal3 10031 -1811 10031 -1811 0 FreeSans 80 0 0 0 SA_OUT[11]
port 300 nsew
flabel metal3 10035 -1890 10035 -1890 0 FreeSans 80 0 0 0 SA_OUT[12]
port 301 nsew
flabel metal3 10031 -1954 10031 -1954 0 FreeSans 80 0 0 0 SA_OUT[13]
port 302 nsew
flabel metal3 10034 -2069 10034 -2069 0 FreeSans 80 0 0 0 SA_OUT[14]
port 303 nsew
flabel metal3 10026 -2158 10026 -2158 0 FreeSans 80 0 0 0 SA_OUT[15]
port 304 nsew
flabel metal3 -4539 -2434 -4539 -2434 0 FreeSans 80 0 0 0 EN
port 305 nsew
flabel metal3 -4536 -2510 -4536 -2510 0 FreeSans 80 0 0 0 PRE_A
port 306 nsew
flabel metal2 -4114 -9024 -4100 -9017 0 FreeSans 80 0 0 0 SAEN
port 180 nsew
flabel metal2 -4048 -9024 -4034 -9017 0 FreeSans 80 0 0 0 VCLP
port 179 nsew
flabel metal2 -3982 -9024 -3968 -9017 0 FreeSans 80 0 0 0 PRE_CLSA
port 178 nsew
flabel metal2 -3136 -9015 -3136 -9015 0 FreeSans 40 0 0 0 ADC0_OUT[0]
port 187 nsew
flabel metal2 -3095 -9008 -3095 -9007 0 FreeSans 40 0 0 0 ADC0_OUT[1]
port 190 nsew
flabel metal2 -3054 -9015 -3054 -9015 0 FreeSans 40 0 0 0 ADC0_OUT[2]
port 191 nsew
flabel metal2 -3014 -9008 -3014 -9008 0 FreeSans 40 0 0 0 ADC0_OUT[3]
port 192 nsew
flabel metal2 -1857 -9000 -1857 -9000 0 FreeSans 40 0 0 0 ADC1_OUT[3]
port 196 nsew
flabel metal2 -1898 -9008 -1898 -9008 0 FreeSans 40 0 0 0 ADC1_OUT[2]
port 195 nsew
flabel metal2 -1940 -9000 -1940 -9000 0 FreeSans 40 0 0 0 ADC1_OUT[1]
port 194 nsew
flabel metal2 -1980 -9007 -1980 -9007 0 FreeSans 40 0 0 0 ADC1_OUT[0]
port 193 nsew
flabel metal2 -812 -8984 -811 -8984 0 FreeSans 40 0 0 0 ADC2_OUT[0]
port 197 nsew
flabel metal2 -771 -8978 -771 -8978 0 FreeSans 40 0 0 0 ADC2_OUT[1]
port 198 nsew
flabel metal2 -729 -8983 -729 -8983 0 FreeSans 40 0 0 0 ADC2_OUT[2]
port 199 nsew
flabel metal2 -688 -8977 -688 -8977 0 FreeSans 40 0 0 0 ADC2_OUT[3]
port 200 nsew
flabel metal2 380 -8976 380 -8976 0 FreeSans 40 0 0 0 ADC3_OUT[0]
port 201 nsew
flabel metal2 420 -8971 420 -8971 0 FreeSans 40 0 0 0 ADC3_OUT[1]
port 202 nsew
flabel metal2 461 -8975 461 -8975 0 FreeSans 40 0 0 0 ADC3_OUT[2]
port 203 nsew
flabel metal2 503 -8968 503 -8968 0 FreeSans 40 0 0 0 ADC3_OUT[3]
port 204 nsew
flabel metal2 1679 -8985 1679 -8985 0 FreeSans 40 0 0 0 ADC4_OUT[3]
port 209 nsew
flabel metal2 1640 -8993 1640 -8993 0 FreeSans 40 0 0 0 ADC4_OUT[2]
port 208 nsew
flabel metal2 1597 -8984 1597 -8984 0 FreeSans 40 0 0 0 ADC4_OUT[1]
port 207 nsew
flabel metal2 1556 -8993 1556 -8993 0 FreeSans 40 0 0 0 ADC4_OUT[0]
port 205 nsew
flabel metal2 2733 -9006 2733 -9006 0 FreeSans 40 0 0 0 ADC5_OUT[0]
port 210 nsew
flabel metal2 2774 -8995 2774 -8995 0 FreeSans 40 0 0 0 ADC5_OUT[1]
port 211 nsew
flabel metal2 2815 -9005 2815 -9005 0 FreeSans 40 0 0 0 ADC5_OUT[2]
port 212 nsew
flabel metal2 2857 -8996 2857 -8996 0 FreeSans 40 0 0 0 ADC5_OUT[3]
port 213 nsew
flabel metal2 3915 -9017 3915 -9017 0 FreeSans 40 0 0 0 ADC6_OUT[0]
port 214 nsew
flabel metal2 3956 -9005 3956 -9005 0 FreeSans 40 0 0 0 ADC6_OUT[1]
port 215 nsew
flabel metal2 3998 -9016 3998 -9016 0 FreeSans 40 0 0 0 ADC6_OUT[2]
port 216 nsew
flabel metal2 4039 -9005 4039 -9005 0 FreeSans 40 0 0 0 ADC6_OUT[3]
port 217 nsew
flabel metal2 5225 -9013 5225 -9013 0 FreeSans 40 0 0 0 ADC7_OUT[3]
port 221 nsew
flabel metal2 5184 -9025 5184 -9025 0 FreeSans 40 0 0 0 ADC7_OUT[2]
port 220 nsew
flabel metal2 5142 -9013 5142 -9013 0 FreeSans 40 0 0 0 ADC7_OUT[1]
port 219 nsew
flabel metal2 5101 -9025 5101 -9025 0 FreeSans 40 0 0 0 ADC7_OUT[0]
port 218 nsew
flabel metal2 6281 -9022 6281 -9022 0 FreeSans 40 0 0 0 ADC8_OUT[0]
port 222 nsew
flabel metal2 6321 -9010 6321 -9010 0 FreeSans 40 0 0 0 ADC8_OUT[1]
port 223 nsew
flabel metal2 6363 -9022 6363 -9022 0 FreeSans 40 0 0 0 ADC8_OUT[2]
port 224 nsew
flabel metal2 6404 -9011 6404 -9011 0 FreeSans 40 0 0 0 ADC8_OUT[3]
port 225 nsew
flabel metal2 7509 -8999 7509 -8999 0 FreeSans 40 0 0 0 ADC9_OUT[1]
port 227 nsew
flabel metal2 7592 -8999 7592 -8999 0 FreeSans 40 0 0 0 ADC9_OUT[3]
port 229 nsew
flabel metal2 7551 -9011 7551 -9011 0 FreeSans 40 0 0 0 ADC9_OUT[2]
port 228 nsew
flabel metal2 7468 -9011 7468 -9011 0 FreeSans 40 0 0 0 ADC9_OUT[0]
port 226 nsew
flabel metal2 8641 -9026 8641 -9026 0 FreeSans 40 0 0 0 ADC10_OUT[0]
port 230 nsew
flabel metal2 8682 -9014 8682 -9014 0 FreeSans 40 0 0 0 ADC10_OUT[1]
port 231 nsew
flabel metal2 8724 -9026 8724 -9026 0 FreeSans 40 0 0 0 ADC10_OUT[2]
port 232 nsew
flabel metal2 8765 -9014 8765 -9014 0 FreeSans 40 0 0 0 ADC10_OUT[3]
port 233 nsew
flabel metal2 9823 -9034 9823 -9034 0 FreeSans 40 0 0 0 ADC11_OUT[0]
port 234 nsew
flabel metal2 9864 -9022 9864 -9022 0 FreeSans 40 0 0 0 ADC11_OUT[1]
port 235 nsew
flabel metal2 9906 -9034 9906 -9034 0 FreeSans 40 0 0 0 ADC11_OUT[2]
port 236 nsew
flabel metal2 9947 -9022 9947 -9022 0 FreeSans 40 0 0 0 ADC11_OUT[3]
port 237 nsew
flabel metal2 11012 -9016 11012 -9016 0 FreeSans 40 0 0 0 ADC12_OUT[0]
port 238 nsew
flabel metal2 11053 -9004 11053 -9004 0 FreeSans 40 0 0 0 ADC12_OUT[1]
port 239 nsew
flabel metal2 11095 -9016 11095 -9016 0 FreeSans 40 0 0 0 ADC12_OUT[2]
port 240 nsew
flabel metal2 11136 -9004 11136 -9004 0 FreeSans 40 0 0 0 ADC12_OUT[3]
port 241 nsew
flabel metal2 12208 -9012 12208 -9012 0 FreeSans 40 0 0 0 ADC13_OUT[0]
port 242 nsew
flabel metal2 12248 -9000 12248 -9000 0 FreeSans 40 0 0 0 ADC13_OUT[1]
port 243 nsew
flabel metal2 12290 -9013 12290 -9013 0 FreeSans 40 0 0 0 ADC13_OUT[2]
port 244 nsew
flabel metal2 12331 -9000 12331 -9000 0 FreeSans 40 0 0 0 ADC13_OUT[3]
port 245 nsew
flabel metal2 13384 -9006 13384 -9006 0 FreeSans 40 0 0 0 ADC14_OUT[0]
port 246 nsew
flabel metal2 13424 -8994 13424 -8994 0 FreeSans 40 0 0 0 ADC14_OUT[1]
port 247 nsew
flabel metal2 13466 -9006 13466 -9006 0 FreeSans 40 0 0 0 ADC14_OUT[2]
port 248 nsew
flabel metal2 13506 -8994 13506 -8994 0 FreeSans 40 0 0 0 ADC14_OUT[3]
port 249 nsew
flabel metal2 14411 -8998 14411 -8998 0 FreeSans 40 0 0 0 ADC15_OUT[3]
port 253 nsew
flabel metal2 14370 -9010 14370 -9010 0 FreeSans 40 0 0 0 ADC15_OUT[2]
port 252 nsew
flabel metal2 14328 -8998 14328 -8998 0 FreeSans 40 0 0 0 ADC15_OUT[1]
port 251 nsew
flabel metal2 14288 -9009 14288 -9009 0 FreeSans 40 0 0 0 ADC15_OUT[0]
port 250 nsew
flabel metal3 -4537 5046 -4537 5046 0 FreeSans 80 0 0 0 VDD
port 307 nsew
flabel metal1 -4549 5000 -4546 5014 0 FreeSans 80 0 0 0 PRE_SRAM
port 85 nsew
flabel metal3 -4541 -2046 -4541 -2046 0 FreeSans 80 0 0 0 VSS
port 308 nsew
flabel metal2 14451 -9009 14468 -9005 0 FreeSans 80 0 0 0 Iref0
port 309 nsew
flabel metal2 14507 -9009 14524 -9005 0 FreeSans 80 0 0 0 Iref1
port 310 nsew
flabel metal2 14561 -9009 14578 -9005 0 FreeSans 80 0 0 0 Iref2
port 311 nsew
flabel metal2 14616 -9009 14633 -9005 0 FreeSans 80 0 0 0 Iref3
port 312 nsew
<< end >>
