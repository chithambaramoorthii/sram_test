VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Integrated_bitcell_with_dummy_cells
  CLASS BLOCK ;
  FOREIGN Integrated_bitcell_with_dummy_cells ;
  ORIGIN 45.520 90.350 ;
  SIZE 191.920 BY 143.910 ;
  PIN PRE_SRAM
    PORT
      LAYER met1 ;
        RECT 92.330 49.960 92.660 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 91.460 49.960 91.790 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.590 49.960 90.920 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.580 49.960 86.910 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 85.710 49.960 86.040 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.840 49.960 85.170 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.830 49.960 81.160 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.960 49.960 80.290 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.090 49.960 79.420 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.080 49.960 75.410 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 74.210 49.960 74.540 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.340 49.960 73.670 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.330 49.960 69.660 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 68.460 49.960 68.790 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.590 49.960 67.920 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.580 49.960 63.910 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 62.710 49.960 63.040 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.840 49.960 62.170 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.830 49.960 58.160 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.960 49.960 57.290 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.090 49.960 56.420 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.080 49.960 52.410 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 51.210 49.960 51.540 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.340 49.960 50.670 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.330 49.960 46.660 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 45.460 49.960 45.790 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.590 49.960 44.920 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.580 49.960 40.910 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 39.710 49.960 40.040 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.840 49.960 39.170 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.830 49.960 35.160 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.960 49.960 34.290 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.090 49.960 33.420 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.080 49.960 29.410 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 28.210 49.960 28.540 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.340 49.960 27.670 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.330 49.960 23.660 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.460 49.960 22.790 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.590 49.960 21.920 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.580 49.960 17.910 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 16.710 49.960 17.040 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.840 49.960 16.170 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.830 49.960 12.160 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.960 49.960 11.290 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.090 49.960 10.420 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.080 49.960 6.410 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.210 49.960 5.540 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.340 49.960 4.670 50.000 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 50.000 94.660 50.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 92.330 50.140 92.660 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 91.460 50.140 91.790 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.590 50.140 90.920 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.580 50.140 86.910 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 85.710 50.140 86.040 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.840 50.140 85.170 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.830 50.140 81.160 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.960 50.140 80.290 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.090 50.140 79.420 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.080 50.140 75.410 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 74.210 50.140 74.540 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.340 50.140 73.670 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.330 50.140 69.660 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 68.460 50.140 68.790 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.590 50.140 67.920 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.580 50.140 63.910 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 62.710 50.140 63.040 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.840 50.140 62.170 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.830 50.140 58.160 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.960 50.140 57.290 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.090 50.140 56.420 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.080 50.140 52.410 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 51.210 50.140 51.540 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.340 50.140 50.670 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.330 50.140 46.660 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 45.460 50.140 45.790 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.590 50.140 44.920 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.580 50.140 40.910 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 39.710 50.140 40.040 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.840 50.140 39.170 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.830 50.140 35.160 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.960 50.140 34.290 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.090 50.140 33.420 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.080 50.140 29.410 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 28.210 50.140 28.540 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.340 50.140 27.670 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.330 50.140 23.660 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.460 50.140 22.790 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.590 50.140 21.920 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.580 50.140 17.910 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 16.710 50.140 17.040 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.840 50.140 16.170 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.830 50.140 12.160 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.960 50.140 11.290 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.090 50.140 10.420 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.080 50.140 6.410 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.210 50.140 5.540 50.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.340 50.140 4.670 50.190 ;
    END
  END PRE_SRAM
  PIN RWL[0]
    PORT
      LAYER met1 ;
        RECT 88.710 37.330 89.010 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 37.330 83.260 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 37.330 77.510 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 37.330 71.760 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 37.330 66.010 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 37.330 60.260 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 37.330 54.510 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 37.330 48.760 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 37.330 43.010 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 37.330 37.260 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 37.330 31.510 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 37.330 25.760 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 37.330 20.010 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 37.330 14.260 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 37.330 8.510 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 37.330 2.760 37.410 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 37.410 94.660 37.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 37.550 89.010 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 37.550 83.260 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 37.550 77.510 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 37.550 71.760 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 37.550 66.010 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 37.550 60.260 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 37.550 54.510 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 37.550 48.760 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 37.550 43.010 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 37.550 37.260 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 37.550 31.510 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 37.550 25.760 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 37.550 20.010 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 37.550 14.260 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 37.550 8.510 37.620 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 37.550 2.760 37.620 ;
    END
  END RWL[0]
  PIN WWL[0]
    PORT
      LAYER met1 ;
        RECT 92.300 36.890 92.590 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 36.890 86.840 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 36.890 81.090 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 36.890 75.340 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 36.890 69.590 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 36.890 63.840 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 36.890 58.090 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 36.890 52.340 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 36.890 46.590 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 36.890 40.840 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 36.890 35.090 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 36.890 29.340 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 36.890 23.590 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 36.890 17.840 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 36.890 12.090 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 36.890 6.340 37.010 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 37.010 94.660 37.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 37.150 90.980 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 37.150 85.230 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 37.150 79.480 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 37.150 73.730 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 37.150 67.980 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 37.150 62.230 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 37.150 56.480 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 37.150 50.730 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 37.150 44.980 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 37.150 39.230 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 37.150 33.480 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 37.150 27.730 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 37.150 21.980 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 37.150 16.230 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 37.150 10.480 37.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 37.150 4.730 37.270 ;
    END
  END WWL[0]
  PIN RWLB[0]
    PORT
      LAYER met1 ;
        RECT 94.260 36.510 94.560 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 36.510 88.810 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 36.510 83.060 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 36.510 77.310 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 36.510 71.560 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 36.510 65.810 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 36.510 60.060 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 36.510 54.310 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 36.510 48.560 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 36.510 42.810 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 36.510 37.060 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 36.510 31.310 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 36.510 25.560 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 36.510 19.810 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 36.510 14.060 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 36.510 8.310 36.600 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 36.600 94.660 36.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 36.740 94.560 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 36.740 88.810 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 36.740 83.060 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 36.740 77.310 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 36.740 71.560 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 36.740 65.810 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 36.740 60.060 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 36.740 54.310 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 36.740 48.560 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 36.740 42.810 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 36.740 37.060 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 36.740 31.310 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 36.740 25.560 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 36.740 19.810 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 36.740 14.060 36.840 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 36.740 8.310 36.840 ;
    END
  END RWLB[0]
  PIN RWL[1]
    PORT
      LAYER met1 ;
        RECT 88.710 34.920 89.010 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 34.920 83.260 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 34.920 77.510 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 34.920 71.760 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 34.920 66.010 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 34.920 60.260 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 34.920 54.510 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 34.920 48.760 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 34.920 43.010 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 34.920 37.260 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 34.920 31.510 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 34.920 25.760 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 34.920 20.010 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 34.920 14.260 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 34.920 8.510 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 34.920 2.760 35.000 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 35.000 94.660 35.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 35.140 89.010 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 35.140 83.260 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 35.140 77.510 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 35.140 71.760 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 35.140 66.010 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 35.140 60.260 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 35.140 54.510 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 35.140 48.760 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 35.140 43.010 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 35.140 37.260 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 35.140 31.510 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 35.140 25.760 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 35.140 20.010 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 35.140 14.260 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 35.140 8.510 35.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 35.140 2.760 35.210 ;
    END
  END RWL[1]
  PIN WWL[1]
    PORT
      LAYER met1 ;
        RECT 92.300 34.480 92.590 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 34.480 86.840 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 34.480 81.090 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 34.480 75.340 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 34.480 69.590 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 34.480 63.840 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 34.480 58.090 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 34.480 52.340 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 34.480 46.590 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 34.480 40.840 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 34.480 35.090 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 34.480 29.340 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 34.480 23.590 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 34.480 17.840 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 34.480 12.090 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 34.480 6.340 34.600 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 34.600 94.660 34.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 34.740 90.980 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 34.740 85.230 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 34.740 79.480 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 34.740 73.730 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 34.740 67.980 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 34.740 62.230 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 34.740 56.480 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 34.740 50.730 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 34.740 44.980 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 34.740 39.230 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 34.740 33.480 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 34.740 27.730 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 34.740 21.980 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 34.740 16.230 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 34.740 10.480 34.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 34.740 4.730 34.860 ;
    END
  END WWL[1]
  PIN RWLB[1]
    PORT
      LAYER met1 ;
        RECT 94.260 34.100 94.560 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 34.100 88.810 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 34.100 83.060 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 34.100 77.310 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 34.100 71.560 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 34.100 65.810 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 34.100 60.060 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 34.100 54.310 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 34.100 48.560 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 34.100 42.810 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 34.100 37.060 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 34.100 31.310 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 34.100 25.560 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 34.100 19.810 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 34.100 14.060 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 34.100 8.310 34.190 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 34.190 94.660 34.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 34.330 94.560 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 34.330 88.810 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 34.330 83.060 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 34.330 77.310 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 34.330 71.560 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 34.330 65.810 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 34.330 60.060 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 34.330 54.310 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 34.330 48.560 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 34.330 42.810 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 34.330 37.060 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 34.330 31.310 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 34.330 25.560 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 34.330 19.810 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 34.330 14.060 34.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 34.330 8.310 34.430 ;
    END
  END RWLB[1]
  PIN RWL[2]
    PORT
      LAYER met1 ;
        RECT 88.710 32.510 89.010 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 32.510 83.260 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 32.510 77.510 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 32.510 71.760 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 32.510 66.010 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 32.510 60.260 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 32.510 54.510 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 32.510 48.760 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 32.510 43.010 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 32.510 37.260 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 32.510 31.510 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 32.510 25.760 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 32.510 20.010 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 32.510 14.260 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 32.510 8.510 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 32.510 2.760 32.590 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 32.590 94.660 32.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 32.730 89.010 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 32.730 83.260 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 32.730 77.510 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 32.730 71.760 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 32.730 66.010 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 32.730 60.260 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 32.730 54.510 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 32.730 48.760 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 32.730 43.010 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 32.730 37.260 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 32.730 31.510 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 32.730 25.760 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 32.730 20.010 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 32.730 14.260 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 32.730 8.510 32.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 32.730 2.760 32.800 ;
    END
  END RWL[2]
  PIN WWL[2]
    PORT
      LAYER met1 ;
        RECT 92.300 32.070 92.590 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 32.070 86.840 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 32.070 81.090 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 32.070 75.340 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 32.070 69.590 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 32.070 63.840 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 32.070 58.090 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 32.070 52.340 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 32.070 46.590 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 32.070 40.840 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 32.070 35.090 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 32.070 29.340 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 32.070 23.590 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 32.070 17.840 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 32.070 12.090 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 32.070 6.340 32.190 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 32.190 94.660 32.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 32.330 90.980 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 32.330 85.230 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 32.330 79.480 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 32.330 73.730 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 32.330 67.980 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 32.330 62.230 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 32.330 56.480 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 32.330 50.730 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 32.330 44.980 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 32.330 39.230 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 32.330 33.480 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 32.330 27.730 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 32.330 21.980 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 32.330 16.230 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 32.330 10.480 32.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 32.330 4.730 32.450 ;
    END
  END WWL[2]
  PIN RWLB[2]
    PORT
      LAYER met1 ;
        RECT 94.260 31.690 94.560 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 31.690 88.810 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 31.690 83.060 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 31.690 77.310 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 31.690 71.560 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 31.690 65.810 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 31.690 60.060 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 31.690 54.310 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 31.690 48.560 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 31.690 42.810 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 31.690 37.060 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 31.690 31.310 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 31.690 25.560 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 31.690 19.810 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 31.690 14.060 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 31.690 8.310 31.780 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 31.780 94.660 31.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 31.920 94.560 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 31.920 88.810 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 31.920 83.060 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 31.920 77.310 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 31.920 71.560 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 31.920 65.810 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 31.920 60.060 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 31.920 54.310 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 31.920 48.560 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 31.920 42.810 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 31.920 37.060 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 31.920 31.310 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 31.920 25.560 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 31.920 19.810 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 31.920 14.060 32.020 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 31.920 8.310 32.020 ;
    END
  END RWLB[2]
  PIN RWL[3]
    PORT
      LAYER met1 ;
        RECT 88.710 30.100 89.010 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 30.100 83.260 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 30.100 77.510 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 30.100 71.760 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 30.100 66.010 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 30.100 60.260 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 30.100 54.510 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 30.100 48.760 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 30.100 43.010 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 30.100 37.260 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 30.100 31.510 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 30.100 25.760 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 30.100 20.010 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 30.100 14.260 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 30.100 8.510 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 30.100 2.760 30.180 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 30.180 94.660 30.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 30.320 89.010 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 30.320 83.260 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 30.320 77.510 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 30.320 71.760 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 30.320 66.010 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 30.320 60.260 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 30.320 54.510 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 30.320 48.760 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 30.320 43.010 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 30.320 37.260 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 30.320 31.510 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 30.320 25.760 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 30.320 20.010 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 30.320 14.260 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 30.320 8.510 30.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 30.320 2.760 30.390 ;
    END
  END RWL[3]
  PIN WWL[3]
    PORT
      LAYER met1 ;
        RECT 92.300 29.660 92.590 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 29.660 86.840 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 29.660 81.090 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 29.660 75.340 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 29.660 69.590 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 29.660 63.840 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 29.660 58.090 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 29.660 52.340 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 29.660 46.590 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 29.660 40.840 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 29.660 35.090 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 29.660 29.340 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 29.660 23.590 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 29.660 17.840 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 29.660 12.090 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 29.660 6.340 29.780 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 29.780 94.660 29.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 29.920 90.980 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 29.920 85.230 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 29.920 79.480 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 29.920 73.730 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 29.920 67.980 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 29.920 62.230 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 29.920 56.480 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 29.920 50.730 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 29.920 44.980 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 29.920 39.230 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 29.920 33.480 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 29.920 27.730 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 29.920 21.980 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 29.920 16.230 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 29.920 10.480 30.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 29.920 4.730 30.040 ;
    END
  END WWL[3]
  PIN RWLB[3]
    PORT
      LAYER met1 ;
        RECT 94.260 29.280 94.560 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 29.280 88.810 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 29.280 83.060 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 29.280 77.310 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 29.280 71.560 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 29.280 65.810 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 29.280 60.060 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 29.280 54.310 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 29.280 48.560 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 29.280 42.810 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 29.280 37.060 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 29.280 31.310 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 29.280 25.560 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 29.280 19.810 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 29.280 14.060 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 29.280 8.310 29.370 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 29.370 94.660 29.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 29.510 94.560 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 29.510 88.810 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 29.510 83.060 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 29.510 77.310 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 29.510 71.560 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 29.510 65.810 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 29.510 60.060 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 29.510 54.310 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 29.510 48.560 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 29.510 42.810 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 29.510 37.060 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 29.510 31.310 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 29.510 25.560 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 29.510 19.810 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 29.510 14.060 29.610 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 29.510 8.310 29.610 ;
    END
  END RWLB[3]
  PIN RWL[4]
    PORT
      LAYER met1 ;
        RECT 88.710 27.290 89.010 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 27.290 83.260 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 27.290 77.510 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 27.290 71.760 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 27.290 66.010 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 27.290 60.260 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 27.290 54.510 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 27.290 48.760 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 27.290 43.010 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 27.290 37.260 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 27.290 31.510 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 27.290 25.760 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 27.290 20.010 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 27.290 14.260 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 27.290 8.510 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 27.290 2.760 27.370 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 27.370 94.660 27.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 27.510 89.010 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 27.510 83.260 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 27.510 77.510 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 27.510 71.760 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 27.510 66.010 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 27.510 60.260 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 27.510 54.510 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 27.510 48.760 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 27.510 43.010 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 27.510 37.260 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 27.510 31.510 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 27.510 25.760 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 27.510 20.010 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 27.510 14.260 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 27.510 8.510 27.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 27.510 2.760 27.570 ;
    END
  END RWL[4]
  PIN WWL[4]
    PORT
      LAYER met1 ;
        RECT 92.300 26.850 92.590 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 26.850 86.840 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 26.850 81.090 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 26.850 75.340 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 26.850 69.590 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 26.850 63.840 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 26.850 58.090 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 26.850 52.340 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 26.850 46.590 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 26.850 40.840 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 26.850 35.090 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 26.850 29.340 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 26.850 23.590 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 26.850 17.840 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 26.850 12.090 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 26.850 6.340 26.970 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 26.970 94.660 27.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 27.110 90.980 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 27.110 85.230 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 27.110 79.480 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 27.110 73.730 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 27.110 67.980 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 27.110 62.230 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 27.110 56.480 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 27.110 50.730 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 27.110 44.980 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 27.110 39.230 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 27.110 33.480 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 27.110 27.730 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 27.110 21.980 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 27.110 16.230 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 27.110 10.480 27.230 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 27.110 4.730 27.230 ;
    END
  END WWL[4]
  PIN RWLB[4]
    PORT
      LAYER met1 ;
        RECT 94.260 26.470 94.560 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 26.470 88.810 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 26.470 83.060 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 26.470 77.310 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 26.470 71.560 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 26.470 65.810 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 26.470 60.060 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 26.470 54.310 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 26.470 48.560 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 26.470 42.810 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 26.470 37.060 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 26.470 31.310 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 26.470 25.560 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 26.470 19.810 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 26.470 14.060 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 26.470 8.310 26.560 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 26.560 94.660 26.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 26.700 94.560 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 26.700 88.810 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 26.700 83.060 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 26.700 77.310 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 26.700 71.560 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 26.700 65.810 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 26.700 60.060 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 26.700 54.310 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 26.700 48.560 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 26.700 42.810 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 26.700 37.060 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 26.700 31.310 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 26.700 25.560 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 26.700 19.810 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 26.700 14.060 26.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 26.700 8.310 26.800 ;
    END
  END RWLB[4]
  PIN RWL[5]
    PORT
      LAYER met1 ;
        RECT 88.710 24.880 89.010 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 24.880 83.260 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 24.880 77.510 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 24.880 71.760 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 24.880 66.010 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 24.880 60.260 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 24.880 54.510 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 24.880 48.760 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 24.880 43.010 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 24.880 37.260 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 24.880 31.510 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 24.880 25.760 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 24.880 20.010 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 24.880 14.260 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 24.880 8.510 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 24.880 2.760 24.960 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 24.960 94.660 25.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 25.100 89.010 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 25.100 83.260 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 25.100 77.510 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 25.100 71.760 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 25.100 66.010 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 25.100 60.260 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 25.100 54.510 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 25.100 48.760 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 25.100 43.010 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 25.100 37.260 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 25.100 31.510 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 25.100 25.760 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 25.100 20.010 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 25.100 14.260 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 25.100 8.510 25.170 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 25.100 2.760 25.170 ;
    END
  END RWL[5]
  PIN WWL[5]
    PORT
      LAYER met1 ;
        RECT 92.300 24.440 92.590 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 24.440 86.840 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 24.440 81.090 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 24.440 75.340 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 24.440 69.590 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 24.440 63.840 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 24.440 58.090 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 24.440 52.340 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 24.440 46.590 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 24.440 40.840 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 24.440 35.090 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 24.440 29.340 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 24.440 23.590 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 24.440 17.840 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 24.440 12.090 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 24.440 6.340 24.560 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 24.560 94.660 24.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 24.700 90.980 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 24.700 85.230 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 24.700 79.480 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 24.700 73.730 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 24.700 67.980 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 24.700 62.230 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 24.700 56.480 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 24.700 50.730 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 24.700 44.980 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 24.700 39.230 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 24.700 33.480 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 24.700 27.730 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 24.700 21.980 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 24.700 16.230 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 24.700 10.480 24.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 24.700 4.730 24.820 ;
    END
  END WWL[5]
  PIN RWLB[5]
    PORT
      LAYER met1 ;
        RECT 94.260 24.060 94.560 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 24.060 88.810 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 24.060 83.060 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 24.060 77.310 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 24.060 71.560 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 24.060 65.810 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 24.060 60.060 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 24.060 54.310 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 24.060 48.560 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 24.060 42.810 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 24.060 37.060 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 24.060 31.310 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 24.060 25.560 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 24.060 19.810 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 24.060 14.060 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 24.060 8.310 24.150 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 24.150 94.660 24.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 24.290 94.560 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 24.290 88.810 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 24.290 83.060 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 24.290 77.310 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 24.290 71.560 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 24.290 65.810 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 24.290 60.060 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 24.290 54.310 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 24.290 48.560 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 24.290 42.810 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 24.290 37.060 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 24.290 31.310 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 24.290 25.560 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 24.290 19.810 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 24.290 14.060 24.390 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 24.290 8.310 24.390 ;
    END
  END RWLB[5]
  PIN RWL[6]
    PORT
      LAYER met1 ;
        RECT 88.710 22.470 89.010 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 22.470 83.260 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 22.470 77.510 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 22.470 71.760 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 22.470 66.010 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 22.470 60.260 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 22.470 54.510 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 22.470 48.760 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 22.470 43.010 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 22.470 37.260 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 22.470 31.510 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 22.470 25.760 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 22.470 20.010 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 22.470 14.260 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 22.470 8.510 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 22.470 2.760 22.550 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 22.550 94.660 22.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 22.690 89.010 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 22.690 83.260 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 22.690 77.510 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 22.690 71.760 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 22.690 66.010 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 22.690 60.260 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 22.690 54.510 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 22.690 48.760 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 22.690 43.010 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 22.690 37.260 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 22.690 31.510 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 22.690 25.760 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 22.690 20.010 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 22.690 14.260 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 22.690 8.510 22.760 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 22.690 2.760 22.760 ;
    END
  END RWL[6]
  PIN WWL[6]
    PORT
      LAYER met1 ;
        RECT 92.300 22.030 92.590 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 22.030 86.840 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 22.030 81.090 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 22.030 75.340 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 22.030 69.590 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 22.030 63.840 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 22.030 58.090 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 22.030 52.340 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 22.030 46.590 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 22.030 40.840 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 22.030 35.090 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 22.030 29.340 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 22.030 23.590 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 22.030 17.840 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 22.030 12.090 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 22.030 6.340 22.150 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 22.150 94.660 22.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 22.290 90.980 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 22.290 85.230 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 22.290 79.480 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 22.290 73.730 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 22.290 67.980 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 22.290 62.230 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 22.290 56.480 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 22.290 50.730 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 22.290 44.980 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 22.290 39.230 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 22.290 33.480 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 22.290 27.730 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 22.290 21.980 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 22.290 16.230 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 22.290 10.480 22.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 22.290 4.730 22.410 ;
    END
  END WWL[6]
  PIN RWLB[6]
    PORT
      LAYER met1 ;
        RECT 94.260 21.650 94.560 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 21.650 88.810 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 21.650 83.060 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 21.650 77.310 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 21.650 71.560 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 21.650 65.810 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 21.650 60.060 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 21.650 54.310 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 21.650 48.560 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 21.650 42.810 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 21.650 37.060 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 21.650 31.310 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 21.650 25.560 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 21.650 19.810 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 21.650 14.060 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 21.650 8.310 21.740 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 21.740 94.660 21.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 21.880 94.560 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 21.880 88.810 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 21.880 83.060 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 21.880 77.310 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 21.880 71.560 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 21.880 65.810 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 21.880 60.060 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 21.880 54.310 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 21.880 48.560 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 21.880 42.810 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 21.880 37.060 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 21.880 31.310 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 21.880 25.560 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 21.880 19.810 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 21.880 14.060 21.980 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 21.880 8.310 21.980 ;
    END
  END RWLB[6]
  PIN RWL[7]
    PORT
      LAYER met1 ;
        RECT 88.710 20.060 89.010 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 20.060 83.260 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 20.060 77.510 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 20.060 71.760 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 20.060 66.010 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 20.060 60.260 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 20.060 54.510 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 20.060 48.760 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 20.060 43.010 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 20.060 37.260 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 20.060 31.510 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 20.060 25.760 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 20.060 20.010 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 20.060 14.260 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 20.060 8.510 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 20.060 2.760 20.140 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 20.140 94.660 20.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 20.280 89.010 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 20.280 83.260 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 20.280 77.510 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 20.280 71.760 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 20.280 66.010 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 20.280 60.260 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 20.280 54.510 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 20.280 48.760 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 20.280 43.010 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 20.280 37.260 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 20.280 31.510 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 20.280 25.760 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 20.280 20.010 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 20.280 14.260 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 20.280 8.510 20.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 20.280 2.760 20.350 ;
    END
  END RWL[7]
  PIN WWL[7]
    PORT
      LAYER met1 ;
        RECT 92.300 19.620 92.590 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 19.620 86.840 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 19.620 81.090 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 19.620 75.340 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 19.620 69.590 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 19.620 63.840 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 19.620 58.090 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 19.620 52.340 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 19.620 46.590 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 19.620 40.840 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 19.620 35.090 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 19.620 29.340 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 19.620 23.590 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 19.620 17.840 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 19.620 12.090 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 19.620 6.340 19.740 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 19.740 94.660 19.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 19.880 90.980 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 19.880 85.230 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 19.880 79.480 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 19.880 73.730 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 19.880 67.980 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 19.880 62.230 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 19.880 56.480 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 19.880 50.730 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 19.880 44.980 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 19.880 39.230 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 19.880 33.480 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 19.880 27.730 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 19.880 21.980 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 19.880 16.230 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 19.880 10.480 20.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 19.880 4.730 20.000 ;
    END
  END WWL[7]
  PIN RWLB[7]
    PORT
      LAYER met1 ;
        RECT 94.260 19.240 94.560 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 19.240 88.810 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 19.240 83.060 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 19.240 77.310 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 19.240 71.560 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 19.240 65.810 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 19.240 60.060 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 19.240 54.310 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 19.240 48.560 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 19.240 42.810 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 19.240 37.060 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 19.240 31.310 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 19.240 25.560 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 19.240 19.810 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 19.240 14.060 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 19.240 8.310 19.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 19.330 94.660 19.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 19.470 94.560 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 19.470 88.810 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 19.470 83.060 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 19.470 77.310 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 19.470 71.560 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 19.470 65.810 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 19.470 60.060 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 19.470 54.310 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 19.470 48.560 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 19.470 42.810 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 19.470 37.060 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 19.470 31.310 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 19.470 25.560 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 19.470 19.810 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 19.470 14.060 19.570 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 19.470 8.310 19.570 ;
    END
  END RWLB[7]
  PIN RWL[8]
    PORT
      LAYER met1 ;
        RECT 88.710 17.650 89.010 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 17.650 83.260 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 17.650 77.510 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 17.650 71.760 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 17.650 66.010 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 17.650 60.260 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 17.650 54.510 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 17.650 48.760 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 17.650 43.010 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 17.650 37.260 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 17.650 31.510 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 17.650 25.760 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 17.650 20.010 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 17.650 14.260 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 17.650 8.510 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 17.650 2.760 17.730 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 17.730 94.660 17.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 17.870 89.010 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 17.870 83.260 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 17.870 77.510 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 17.870 71.760 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 17.870 66.010 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 17.870 60.260 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 17.870 54.510 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 17.870 48.760 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 17.870 43.010 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 17.870 37.260 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 17.870 31.510 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 17.870 25.760 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 17.870 20.010 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 17.870 14.260 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 17.870 8.510 17.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 17.870 2.760 17.940 ;
    END
  END RWL[8]
  PIN WWL[8]
    PORT
      LAYER met1 ;
        RECT 92.300 17.210 92.590 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 17.210 86.840 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 17.210 81.090 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 17.210 75.340 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 17.210 69.590 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 17.210 63.840 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 17.210 58.090 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 17.210 52.340 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 17.210 46.590 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 17.210 40.840 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 17.210 35.090 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 17.210 29.340 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 17.210 23.590 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 17.210 17.840 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 17.210 12.090 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 17.210 6.340 17.330 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 17.330 94.660 17.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 17.470 90.980 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 17.470 85.230 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 17.470 79.480 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 17.470 73.730 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 17.470 67.980 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 17.470 62.230 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 17.470 56.480 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 17.470 50.730 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 17.470 44.980 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 17.470 39.230 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 17.470 33.480 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 17.470 27.730 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 17.470 21.980 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 17.470 16.230 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 17.470 10.480 17.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 17.470 4.730 17.590 ;
    END
  END WWL[8]
  PIN RWLB[8]
    PORT
      LAYER met1 ;
        RECT 94.260 16.830 94.560 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 16.830 88.810 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 16.830 83.060 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 16.830 77.310 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 16.830 71.560 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 16.830 65.810 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 16.830 60.060 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 16.830 54.310 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 16.830 48.560 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 16.830 42.810 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 16.830 37.060 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 16.830 31.310 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 16.830 25.560 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 16.830 19.810 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 16.830 14.060 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 16.830 8.310 16.920 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 16.920 94.660 17.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 17.060 94.560 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 17.060 88.810 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 17.060 83.060 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 17.060 77.310 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 17.060 71.560 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 17.060 65.810 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 17.060 60.060 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 17.060 54.310 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 17.060 48.560 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 17.060 42.810 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 17.060 37.060 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 17.060 31.310 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 17.060 25.560 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 17.060 19.810 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 17.060 14.060 17.160 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 17.060 8.310 17.160 ;
    END
  END RWLB[8]
  PIN RWL[9]
    PORT
      LAYER met1 ;
        RECT 88.710 15.240 89.010 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 15.240 83.260 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 15.240 77.510 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 15.240 71.760 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 15.240 66.010 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 15.240 60.260 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 15.240 54.510 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 15.240 48.760 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 15.240 43.010 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 15.240 37.260 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 15.240 31.510 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 15.240 25.760 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 15.240 20.010 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 15.240 14.260 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 15.240 8.510 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 15.240 2.760 15.320 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 15.320 94.660 15.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 15.460 89.010 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 15.460 83.260 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 15.460 77.510 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 15.460 71.760 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 15.460 66.010 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 15.460 60.260 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 15.460 54.510 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 15.460 48.760 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 15.460 43.010 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 15.460 37.260 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 15.460 31.510 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 15.460 25.760 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 15.460 20.010 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 15.460 14.260 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 15.460 8.510 15.530 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 15.460 2.760 15.530 ;
    END
  END RWL[9]
  PIN WWL[9]
    PORT
      LAYER met1 ;
        RECT 92.300 14.800 92.590 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 14.800 86.840 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 14.800 81.090 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 14.800 75.340 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 14.800 69.590 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 14.800 63.840 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 14.800 58.090 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 14.800 52.340 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 14.800 46.590 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 14.800 40.840 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 14.800 35.090 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 14.800 29.340 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 14.800 23.590 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 14.800 17.840 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 14.800 12.090 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 14.800 6.340 14.920 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 14.920 94.660 15.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 15.060 90.980 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 15.060 85.230 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 15.060 79.480 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 15.060 73.730 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 15.060 67.980 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 15.060 62.230 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 15.060 56.480 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 15.060 50.730 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 15.060 44.980 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 15.060 39.230 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 15.060 33.480 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 15.060 27.730 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 15.060 21.980 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 15.060 16.230 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 15.060 10.480 15.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 15.060 4.730 15.180 ;
    END
  END WWL[9]
  PIN RWLB[9]
    PORT
      LAYER met1 ;
        RECT 94.260 14.420 94.560 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 14.420 88.810 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 14.420 83.060 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 14.420 77.310 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 14.420 71.560 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 14.420 65.810 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 14.420 60.060 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 14.420 54.310 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 14.420 48.560 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 14.420 42.810 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 14.420 37.060 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 14.420 31.310 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 14.420 25.560 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 14.420 19.810 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 14.420 14.060 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 14.420 8.310 14.510 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 14.510 94.660 14.650 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 14.650 94.560 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 14.650 88.810 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 14.650 83.060 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 14.650 77.310 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 14.650 71.560 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 14.650 65.810 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 14.650 60.060 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 14.650 54.310 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 14.650 48.560 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 14.650 42.810 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 14.650 37.060 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 14.650 31.310 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 14.650 25.560 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 14.650 19.810 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 14.650 14.060 14.750 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 14.650 8.310 14.750 ;
    END
  END RWLB[9]
  PIN RWL[10]
    PORT
      LAYER met1 ;
        RECT 88.710 12.830 89.010 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 12.830 83.260 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 12.830 77.510 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 12.830 71.760 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 12.830 66.010 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 12.830 60.260 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 12.830 54.510 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 12.830 48.760 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 12.830 43.010 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 12.830 37.260 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 12.830 31.510 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 12.830 25.760 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 12.830 20.010 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 12.830 14.260 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 12.830 8.510 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 12.830 2.760 12.910 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 12.910 94.660 13.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 13.050 89.010 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 13.050 83.260 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 13.050 77.510 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 13.050 71.760 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 13.050 66.010 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 13.050 60.260 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 13.050 54.510 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 13.050 48.760 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 13.050 43.010 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 13.050 37.260 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 13.050 31.510 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 13.050 25.760 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 13.050 20.010 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 13.050 14.260 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 13.050 8.510 13.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 13.050 2.760 13.120 ;
    END
  END RWL[10]
  PIN WWL[10]
    PORT
      LAYER met1 ;
        RECT 92.300 12.390 92.590 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 12.390 86.840 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 12.390 81.090 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 12.390 75.340 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 12.390 69.590 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 12.390 63.840 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 12.390 58.090 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 12.390 52.340 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 12.390 46.590 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 12.390 40.840 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 12.390 35.090 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 12.390 29.340 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 12.390 23.590 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 12.390 17.840 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 12.390 12.090 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 12.390 6.340 12.510 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 12.510 94.660 12.650 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 12.650 90.980 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 12.650 85.230 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 12.650 79.480 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 12.650 73.730 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 12.650 67.980 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 12.650 62.230 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 12.650 56.480 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 12.650 50.730 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 12.650 44.980 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 12.650 39.230 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 12.650 33.480 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 12.650 27.730 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 12.650 21.980 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 12.650 16.230 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 12.650 10.480 12.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 12.650 4.730 12.770 ;
    END
  END WWL[10]
  PIN RWLB[10]
    PORT
      LAYER met1 ;
        RECT 94.260 12.010 94.560 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 12.010 88.810 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 12.010 83.060 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 12.010 77.310 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 12.010 71.560 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 12.010 65.810 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 12.010 60.060 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 12.010 54.310 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 12.010 48.560 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 12.010 42.810 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 12.010 37.060 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 12.010 31.310 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 12.010 25.560 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 12.010 19.810 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 12.010 14.060 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 12.010 8.310 12.100 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 12.100 94.660 12.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 12.240 94.560 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 12.240 88.810 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 12.240 83.060 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 12.240 77.310 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 12.240 71.560 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 12.240 65.810 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 12.240 60.060 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 12.240 54.310 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 12.240 48.560 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 12.240 42.810 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 12.240 37.060 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 12.240 31.310 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 12.240 25.560 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 12.240 19.810 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 12.240 14.060 12.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 12.240 8.310 12.340 ;
    END
  END RWLB[10]
  PIN RWL[11]
    PORT
      LAYER met1 ;
        RECT 88.710 10.420 89.010 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 10.420 83.260 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 10.420 77.510 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 10.420 71.760 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 10.420 66.010 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 10.420 60.260 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 10.420 54.510 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 10.420 48.760 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 10.420 43.010 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 10.420 37.260 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 10.420 31.510 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 10.420 25.760 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 10.420 20.010 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 10.420 14.260 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 10.420 8.510 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 10.420 2.760 10.500 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 10.500 94.660 10.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 10.640 89.010 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 10.640 83.260 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 10.640 77.510 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 10.640 71.760 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 10.640 66.010 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 10.640 60.260 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 10.640 54.510 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 10.640 48.760 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 10.640 43.010 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 10.640 37.260 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 10.640 31.510 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 10.640 25.760 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 10.640 20.010 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 10.640 14.260 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 10.640 8.510 10.710 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 10.640 2.760 10.710 ;
    END
  END RWL[11]
  PIN WWL[11]
    PORT
      LAYER met1 ;
        RECT 92.300 9.980 92.590 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 9.980 86.840 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 9.980 81.090 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 9.980 75.340 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 9.980 69.590 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 9.980 63.840 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 9.980 58.090 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 9.980 52.340 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 9.980 46.590 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 9.980 40.840 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 9.980 35.090 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 9.980 29.340 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 9.980 23.590 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 9.980 17.840 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 9.980 12.090 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 9.980 6.340 10.100 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 10.100 94.660 10.240 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 10.240 90.980 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 10.240 85.230 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 10.240 79.480 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 10.240 73.730 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 10.240 67.980 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 10.240 62.230 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 10.240 56.480 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 10.240 50.730 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 10.240 44.980 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 10.240 39.230 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 10.240 33.480 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 10.240 27.730 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 10.240 21.980 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 10.240 16.230 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 10.240 10.480 10.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 10.240 4.730 10.360 ;
    END
  END WWL[11]
  PIN RWLB[11]
    PORT
      LAYER met1 ;
        RECT 94.260 9.600 94.560 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 9.600 88.810 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 9.600 83.060 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 9.600 77.310 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 9.600 71.560 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 9.600 65.810 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 9.600 60.060 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 9.600 54.310 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 9.600 48.560 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 9.600 42.810 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 9.600 37.060 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 9.600 31.310 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 9.600 25.560 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 9.600 19.810 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 9.600 14.060 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 9.600 8.310 9.690 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 9.690 94.660 9.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 9.830 94.560 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 9.830 88.810 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 9.830 83.060 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 9.830 77.310 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 9.830 71.560 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 9.830 65.810 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 9.830 60.060 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 9.830 54.310 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 9.830 48.560 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 9.830 42.810 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 9.830 37.060 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 9.830 31.310 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 9.830 25.560 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 9.830 19.810 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 9.830 14.060 9.930 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 9.830 8.310 9.930 ;
    END
  END RWLB[11]
  PIN RWL[12]
    PORT
      LAYER met1 ;
        RECT 88.710 7.600 89.010 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 7.600 83.260 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 7.600 77.510 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 7.600 71.760 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 7.600 66.010 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 7.600 60.260 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 7.600 54.510 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 7.600 48.760 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 7.600 43.010 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 7.600 37.260 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 7.600 31.510 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 7.600 25.760 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 7.600 20.010 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 7.600 14.260 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 7.600 8.510 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 7.600 2.760 7.680 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 7.680 94.660 7.820 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 7.820 89.010 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 7.820 83.260 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 7.820 77.510 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 7.820 71.760 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 7.820 66.010 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 7.820 60.260 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 7.820 54.510 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 7.820 48.760 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 7.820 43.010 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 7.820 37.260 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 7.820 31.510 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 7.820 25.760 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 7.820 20.010 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 7.820 14.260 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 7.820 8.510 7.880 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 7.820 2.760 7.880 ;
    END
  END RWL[12]
  PIN WWL[12]
    PORT
      LAYER met1 ;
        RECT 92.300 7.160 92.590 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 7.160 86.840 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 7.160 81.090 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 7.160 75.340 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 7.160 69.590 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 7.160 63.840 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 7.160 58.090 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 7.160 52.340 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 7.160 46.590 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 7.160 40.840 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 7.160 35.090 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 7.160 29.340 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 7.160 23.590 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 7.160 17.840 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 7.160 12.090 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 7.160 6.340 7.280 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 7.280 94.660 7.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 7.420 90.980 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 7.420 85.230 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 7.420 79.480 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 7.420 73.730 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 7.420 67.980 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 7.420 62.230 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 7.420 56.480 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 7.420 50.730 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 7.420 44.980 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 7.420 39.230 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 7.420 33.480 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 7.420 27.730 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 7.420 21.980 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 7.420 16.230 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 7.420 10.480 7.540 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 7.420 4.730 7.540 ;
    END
  END WWL[12]
  PIN RWLB[12]
    PORT
      LAYER met1 ;
        RECT 94.260 6.780 94.560 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 6.780 88.810 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 6.780 83.060 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 6.780 77.310 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 6.780 71.560 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 6.780 65.810 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 6.780 60.060 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 6.780 54.310 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 6.780 48.560 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 6.780 42.810 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 6.780 37.060 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 6.780 31.310 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 6.780 25.560 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 6.780 19.810 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 6.780 14.060 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 6.780 8.310 6.870 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 6.870 94.660 7.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 7.010 94.560 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 7.010 88.810 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 7.010 83.060 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 7.010 77.310 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 7.010 71.560 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 7.010 65.810 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 7.010 60.060 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 7.010 54.310 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 7.010 48.560 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 7.010 42.810 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 7.010 37.060 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 7.010 31.310 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 7.010 25.560 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 7.010 19.810 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 7.010 14.060 7.110 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 7.010 8.310 7.110 ;
    END
  END RWLB[12]
  PIN RWL[13]
    PORT
      LAYER met1 ;
        RECT 88.710 5.190 89.010 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 5.190 83.260 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 5.190 77.510 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 5.190 71.760 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 5.190 66.010 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 5.190 60.260 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 5.190 54.510 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 5.190 48.760 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 5.190 43.010 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 5.190 37.260 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 5.190 31.510 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 5.190 25.760 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 5.190 20.010 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 5.190 14.260 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 5.190 8.510 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 5.190 2.760 5.270 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 5.270 94.660 5.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 5.410 89.010 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 5.410 83.260 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 5.410 77.510 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 5.410 71.760 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 5.410 66.010 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 5.410 60.260 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 5.410 54.510 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 5.410 48.760 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 5.410 43.010 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 5.410 37.260 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 5.410 31.510 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 5.410 25.760 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 5.410 20.010 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 5.410 14.260 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 5.410 8.510 5.480 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 5.410 2.760 5.480 ;
    END
  END RWL[13]
  PIN WWL[13]
    PORT
      LAYER met1 ;
        RECT 92.300 4.750 92.590 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 4.750 86.840 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 4.750 81.090 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 4.750 75.340 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 4.750 69.590 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 4.750 63.840 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 4.750 58.090 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 4.750 52.340 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 4.750 46.590 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 4.750 40.840 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 4.750 35.090 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 4.750 29.340 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 4.750 23.590 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 4.750 17.840 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 4.750 12.090 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 4.750 6.340 4.870 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 4.870 94.660 5.010 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 5.010 90.980 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 5.010 85.230 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 5.010 79.480 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 5.010 73.730 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 5.010 67.980 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 5.010 62.230 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 5.010 56.480 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 5.010 50.730 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 5.010 44.980 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 5.010 39.230 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 5.010 33.480 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 5.010 27.730 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 5.010 21.980 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 5.010 16.230 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 5.010 10.480 5.130 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 5.010 4.730 5.130 ;
    END
  END WWL[13]
  PIN RWLB[13]
    PORT
      LAYER met1 ;
        RECT 94.260 4.370 94.560 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 4.370 88.810 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 4.370 83.060 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 4.370 77.310 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 4.370 71.560 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 4.370 65.810 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 4.370 60.060 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 4.370 54.310 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 4.370 48.560 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 4.370 42.810 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 4.370 37.060 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 4.370 31.310 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 4.370 25.560 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 4.370 19.810 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 4.370 14.060 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 4.370 8.310 4.460 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 4.460 94.660 4.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 4.600 94.560 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 4.600 88.810 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 4.600 83.060 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 4.600 77.310 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 4.600 71.560 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 4.600 65.810 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 4.600 60.060 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 4.600 54.310 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 4.600 48.560 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 4.600 42.810 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 4.600 37.060 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 4.600 31.310 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 4.600 25.560 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 4.600 19.810 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 4.600 14.060 4.700 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 4.600 8.310 4.700 ;
    END
  END RWLB[13]
  PIN RWL[14]
    PORT
      LAYER met1 ;
        RECT 88.710 2.780 89.010 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 2.780 83.260 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 2.780 77.510 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 2.780 71.760 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 2.780 66.010 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 2.780 60.260 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 2.780 54.510 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 2.780 48.760 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 2.780 43.010 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 2.780 37.260 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 2.780 31.510 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 2.780 25.760 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 2.780 20.010 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 2.780 14.260 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 2.780 8.510 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 2.780 2.760 2.860 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 2.860 94.660 3.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 3.000 89.010 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 3.000 83.260 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 3.000 77.510 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 3.000 71.760 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 3.000 66.010 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 3.000 60.260 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 3.000 54.510 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 3.000 48.760 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 3.000 43.010 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 3.000 37.260 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 3.000 31.510 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 3.000 25.760 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 3.000 20.010 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 3.000 14.260 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 3.000 8.510 3.070 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 3.000 2.760 3.070 ;
    END
  END RWL[14]
  PIN WWL[14]
    PORT
      LAYER met1 ;
        RECT 92.300 2.340 92.590 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 2.340 86.840 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 2.340 81.090 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 2.340 75.340 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 2.340 69.590 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 2.340 63.840 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 2.340 58.090 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 2.340 52.340 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 2.340 46.590 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 2.340 40.840 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 2.340 35.090 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 2.340 29.340 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 2.340 23.590 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 2.340 17.840 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 2.340 12.090 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 2.340 6.340 2.460 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 2.460 94.660 2.600 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 2.600 90.980 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 2.600 85.230 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 2.600 79.480 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 2.600 73.730 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 2.600 67.980 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 2.600 62.230 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 2.600 56.480 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 2.600 50.730 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 2.600 44.980 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 2.600 39.230 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 2.600 33.480 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 2.600 27.730 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 2.600 21.980 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 2.600 16.230 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 2.600 10.480 2.720 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 2.600 4.730 2.720 ;
    END
  END WWL[14]
  PIN RWLB[14]
    PORT
      LAYER met1 ;
        RECT 94.260 1.960 94.560 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 1.960 88.810 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 1.960 83.060 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 1.960 77.310 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 1.960 71.560 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 1.960 65.810 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 1.960 60.060 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 1.960 54.310 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 1.960 48.560 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 1.960 42.810 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 1.960 37.060 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 1.960 31.310 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 1.960 25.560 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 1.960 19.810 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 1.960 14.060 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 1.960 8.310 2.050 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 2.050 94.660 2.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 2.190 94.560 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 2.190 88.810 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 2.190 83.060 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 2.190 77.310 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 2.190 71.560 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 2.190 65.810 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 2.190 60.060 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 2.190 54.310 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 2.190 48.560 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 2.190 42.810 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 2.190 37.060 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 2.190 31.310 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 2.190 25.560 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 2.190 19.810 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 2.190 14.060 2.290 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 2.190 8.310 2.290 ;
    END
  END RWLB[14]
  PIN RWL[15]
    PORT
      LAYER met1 ;
        RECT 88.710 0.370 89.010 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 0.370 83.260 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 0.370 77.510 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 0.370 71.760 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 0.370 66.010 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 0.370 60.260 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 0.370 54.510 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 0.370 48.760 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 0.370 43.010 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 0.370 37.260 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 0.370 31.510 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 0.370 25.760 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 0.370 20.010 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 0.370 14.260 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 0.370 8.510 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 0.370 2.760 0.450 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 0.450 94.660 0.590 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.710 0.590 89.010 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.960 0.590 83.260 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.210 0.590 77.510 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.460 0.590 71.760 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.710 0.590 66.010 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.960 0.590 60.260 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.210 0.590 54.510 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.460 0.590 48.760 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.710 0.590 43.010 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.960 0.590 37.260 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.210 0.590 31.510 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.460 0.590 25.760 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.710 0.590 20.010 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.960 0.590 14.260 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.210 0.590 8.510 0.660 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.460 0.590 2.760 0.660 ;
    END
  END RWL[15]
  PIN WWL[15]
    PORT
      LAYER met1 ;
        RECT 92.300 -0.070 92.590 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 -0.070 86.840 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 -0.070 81.090 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 -0.070 75.340 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 -0.070 69.590 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 -0.070 63.840 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 -0.070 58.090 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 -0.070 52.340 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 -0.070 46.590 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 -0.070 40.840 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 -0.070 35.090 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 -0.070 29.340 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 -0.070 23.590 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 -0.070 17.840 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 -0.070 12.090 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 -0.070 6.340 0.050 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 0.050 94.660 0.190 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 0.190 90.980 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 0.190 85.230 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 0.190 79.480 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 0.190 73.730 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 0.190 67.980 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 0.190 62.230 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 0.190 56.480 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 0.190 50.730 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 0.190 44.980 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 0.190 39.230 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 0.190 33.480 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 0.190 27.730 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 0.190 21.980 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 0.190 16.230 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 0.190 10.480 0.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 0.190 4.730 0.310 ;
    END
  END WWL[15]
  PIN RWLB[15]
    PORT
      LAYER met1 ;
        RECT 94.260 -0.450 94.560 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 -0.450 88.810 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 -0.450 83.060 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 -0.450 77.310 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 -0.450 71.560 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 -0.450 65.810 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 -0.450 60.060 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 -0.450 54.310 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 -0.450 48.560 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 -0.450 42.810 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 -0.450 37.060 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 -0.450 31.310 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 -0.450 25.560 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 -0.450 19.810 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 -0.450 14.060 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 -0.450 8.310 -0.360 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 -0.360 94.660 -0.220 ;
    END
    PORT
      LAYER met1 ;
        RECT 94.260 -0.220 94.560 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 88.510 -0.220 88.810 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 82.760 -0.220 83.060 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 77.010 -0.220 77.310 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 71.260 -0.220 71.560 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 65.510 -0.220 65.810 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.760 -0.220 60.060 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 54.010 -0.220 54.310 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.260 -0.220 48.560 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 42.510 -0.220 42.810 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 36.760 -0.220 37.060 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 31.010 -0.220 31.310 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 25.260 -0.220 25.560 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 19.510 -0.220 19.810 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 13.760 -0.220 14.060 -0.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 8.010 -0.220 8.310 -0.120 ;
    END
  END RWLB[15]
  PIN PRE_VLSA
    PORT
      LAYER met2 ;
        RECT 93.330 -18.780 93.660 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 93.470 -18.450 93.610 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 89.650 -18.770 89.980 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 87.580 -18.780 87.910 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 89.670 -18.440 89.810 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 87.720 -18.450 87.860 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 83.900 -18.770 84.230 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 81.830 -18.780 82.160 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 83.920 -18.440 84.060 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 81.970 -18.450 82.110 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 78.150 -18.770 78.480 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 76.080 -18.780 76.410 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 78.170 -18.440 78.310 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 76.220 -18.450 76.360 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 72.400 -18.770 72.730 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 70.330 -18.780 70.660 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 72.420 -18.440 72.560 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 70.470 -18.450 70.610 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 66.650 -18.770 66.980 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 64.580 -18.780 64.910 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 66.670 -18.440 66.810 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 64.720 -18.450 64.860 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 60.900 -18.770 61.230 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 58.830 -18.780 59.160 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 60.920 -18.440 61.060 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 58.970 -18.450 59.110 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 55.150 -18.770 55.480 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 53.080 -18.780 53.410 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 55.170 -18.440 55.310 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 53.220 -18.450 53.360 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 49.400 -18.770 49.730 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 47.330 -18.780 47.660 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 49.420 -18.440 49.560 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 47.470 -18.450 47.610 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 43.650 -18.770 43.980 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 41.580 -18.780 41.910 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 43.670 -18.440 43.810 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 41.720 -18.450 41.860 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 37.900 -18.770 38.230 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 35.830 -18.780 36.160 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 37.920 -18.440 38.060 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 35.970 -18.450 36.110 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.150 -18.770 32.480 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.080 -18.780 30.410 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.170 -18.440 32.310 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.220 -18.450 30.360 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 26.400 -18.770 26.730 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 24.330 -18.780 24.660 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 26.420 -18.440 26.560 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 24.470 -18.450 24.610 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 20.650 -18.770 20.980 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 18.580 -18.780 18.910 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 20.670 -18.440 20.810 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 18.720 -18.450 18.860 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.900 -18.770 15.230 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 12.830 -18.780 13.160 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.920 -18.440 15.060 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 12.970 -18.450 13.110 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.150 -18.770 9.480 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.080 -18.780 7.410 -18.450 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.170 -18.440 9.310 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.220 -18.450 7.360 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.400 -18.770 3.730 -18.440 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.420 -18.440 3.560 -14.570 ;
    END
    PORT
      LAYER met2 ;
        RECT 93.370 -14.570 93.690 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 89.580 -14.570 89.910 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 87.620 -14.570 87.940 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 83.830 -14.570 84.160 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 81.870 -14.570 82.190 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 78.080 -14.570 78.410 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 76.120 -14.570 76.440 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 72.330 -14.570 72.660 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 70.370 -14.570 70.690 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 66.580 -14.570 66.910 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 64.620 -14.570 64.940 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 60.830 -14.570 61.160 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 58.870 -14.570 59.190 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 55.080 -14.570 55.410 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 53.120 -14.570 53.440 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 49.330 -14.570 49.660 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 47.370 -14.570 47.690 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 43.580 -14.570 43.910 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 41.620 -14.570 41.940 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 37.830 -14.570 38.160 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 35.870 -14.570 36.190 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.080 -14.570 32.410 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 30.120 -14.570 30.440 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 26.330 -14.570 26.660 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 24.370 -14.570 24.690 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 20.580 -14.570 20.910 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 18.620 -14.570 18.940 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 14.830 -14.570 15.160 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 12.870 -14.570 13.190 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 9.080 -14.570 9.410 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 7.120 -14.570 7.440 -14.240 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.330 -14.570 3.660 -14.240 ;
    END
  END PRE_VLSA
  PIN WE
    PORT
      LAYER met1 ;
        RECT 92.400 -19.690 92.730 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.520 -19.690 90.850 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.650 -19.690 86.980 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.770 -19.690 85.100 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.900 -19.690 81.230 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.020 -19.690 79.350 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.150 -19.690 75.480 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.270 -19.690 73.600 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.400 -19.690 69.730 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.520 -19.690 67.850 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.650 -19.690 63.980 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.770 -19.690 62.100 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.900 -19.690 58.230 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.020 -19.690 56.350 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.150 -19.690 52.480 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.270 -19.690 50.600 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.400 -19.690 46.730 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.520 -19.690 44.850 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.650 -19.690 40.980 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.770 -19.690 39.100 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.900 -19.690 35.230 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.020 -19.690 33.350 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.150 -19.690 29.480 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.270 -19.690 27.600 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.400 -19.690 23.730 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.520 -19.690 21.850 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.650 -19.690 17.980 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.770 -19.690 16.100 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.900 -19.690 12.230 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.020 -19.690 10.350 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.150 -19.690 6.480 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.270 -19.690 4.600 -19.640 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 -19.640 94.660 -19.500 ;
    END
    PORT
      LAYER met1 ;
        RECT 92.400 -19.500 92.730 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.520 -19.500 90.850 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.650 -19.500 86.980 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.770 -19.500 85.100 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.900 -19.500 81.230 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.020 -19.500 79.350 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.150 -19.500 75.480 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.270 -19.500 73.600 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.400 -19.500 69.730 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.520 -19.500 67.850 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.650 -19.500 63.980 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.770 -19.500 62.100 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.900 -19.500 58.230 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.020 -19.500 56.350 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.150 -19.500 52.480 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.270 -19.500 50.600 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.400 -19.500 46.730 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.520 -19.500 44.850 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.650 -19.500 40.980 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.770 -19.500 39.100 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.900 -19.500 35.230 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.020 -19.500 33.350 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.150 -19.500 29.480 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.270 -19.500 27.600 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.400 -19.500 23.730 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.520 -19.500 21.850 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.650 -19.500 17.980 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.770 -19.500 16.100 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.900 -19.500 12.230 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.020 -19.500 10.350 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.150 -19.500 6.480 -19.440 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.270 -19.500 4.600 -19.440 ;
    END
  END WE
  PIN PRE_CLSA
    PORT
      LAYER met2 ;
        RECT -39.820 -90.250 -39.680 -86.190 ;
    END
    PORT
      LAYER met2 ;
        RECT -39.910 -86.190 -39.590 -85.870 ;
    END
    PORT
      LAYER met2 ;
        RECT -39.820 -85.870 -39.680 -58.860 ;
    END
    PORT
      LAYER met2 ;
        RECT -39.870 -58.860 -39.610 -58.540 ;
    END
    PORT
      LAYER met2 ;
        RECT -39.820 -58.540 -39.680 -31.540 ;
    END
    PORT
      LAYER met2 ;
        RECT -39.880 -31.540 -39.620 -31.220 ;
    END
  END PRE_CLSA
  PIN VCLP
    PORT
      LAYER met2 ;
        RECT -40.480 -90.250 -40.340 -81.160 ;
    END
    PORT
      LAYER met2 ;
        RECT -40.570 -81.160 -40.250 -80.840 ;
    END
    PORT
      LAYER met2 ;
        RECT -40.480 -80.840 -40.340 -63.900 ;
    END
    PORT
      LAYER met2 ;
        RECT -40.570 -63.900 -40.250 -63.580 ;
    END
    PORT
      LAYER met2 ;
        RECT -40.480 -63.580 -40.340 -53.830 ;
    END
    PORT
      LAYER met2 ;
        RECT -40.540 -53.830 -40.280 -53.510 ;
    END
    PORT
      LAYER met2 ;
        RECT -40.480 -53.510 -40.340 -36.570 ;
    END
    PORT
      LAYER met2 ;
        RECT -40.540 -36.570 -40.280 -36.250 ;
    END
  END VCLP
  PIN SAEN
    PORT
      LAYER met2 ;
        RECT -41.140 -90.250 -41.000 -80.760 ;
    END
    PORT
      LAYER met2 ;
        RECT -41.230 -80.760 -40.910 -80.440 ;
    END
    PORT
      LAYER met2 ;
        RECT -41.140 -80.440 -41.000 -64.300 ;
    END
    PORT
      LAYER met2 ;
        RECT -41.230 -64.300 -40.910 -63.980 ;
    END
    PORT
      LAYER met2 ;
        RECT -41.140 -63.980 -41.000 -53.430 ;
    END
    PORT
      LAYER met2 ;
        RECT -41.230 -53.430 -40.910 -53.110 ;
    END
    PORT
      LAYER met2 ;
        RECT -41.140 -53.110 -41.000 -36.970 ;
    END
    PORT
      LAYER met2 ;
        RECT -41.200 -36.970 -40.940 -36.650 ;
    END
  END SAEN
  PIN ADC0_OUT[0]
    PORT
      LAYER met2 ;
        RECT -31.420 -90.170 -31.280 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT -31.480 -36.130 -31.220 -35.810 ;
    END
  END ADC0_OUT[0]
  PIN ADC0_OUT[1]
    PORT
      LAYER met2 ;
        RECT -31.010 -90.170 -30.870 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT -31.070 -54.260 -30.810 -53.940 ;
    END
  END ADC0_OUT[1]
  PIN ADC0_OUT[2]
    PORT
      LAYER met2 ;
        RECT -30.610 -90.170 -30.470 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT -30.670 -63.460 -30.410 -63.140 ;
    END
  END ADC0_OUT[2]
  PIN ADC0_OUT[3]
    PORT
      LAYER met2 ;
        RECT -30.200 -90.170 -30.060 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT -30.260 -81.590 -30.000 -81.270 ;
    END
  END ADC0_OUT[3]
  PIN ADC1_OUT[0]
    PORT
      LAYER met2 ;
        RECT -19.870 -90.090 -19.730 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT -19.930 -36.130 -19.670 -35.810 ;
    END
  END ADC1_OUT[0]
  PIN ADC1_OUT[1]
    PORT
      LAYER met2 ;
        RECT -19.470 -90.090 -19.330 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT -19.530 -54.260 -19.270 -53.940 ;
    END
  END ADC1_OUT[1]
  PIN ADC1_OUT[2]
    PORT
      LAYER met2 ;
        RECT -19.050 -90.090 -18.910 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT -19.140 -63.460 -18.820 -63.140 ;
    END
  END ADC1_OUT[2]
  PIN ADC1_OUT[3]
    PORT
      LAYER met2 ;
        RECT -18.640 -90.090 -18.500 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT -18.700 -81.590 -18.440 -81.270 ;
    END
  END ADC1_OUT[3]
  PIN ADC2_OUT[0]
    PORT
      LAYER met2 ;
        RECT -8.180 -89.860 -8.040 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT -8.240 -36.130 -7.980 -35.810 ;
    END
  END ADC2_OUT[0]
  PIN ADC2_OUT[1]
    PORT
      LAYER met2 ;
        RECT -7.780 -89.860 -7.640 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT -7.840 -54.260 -7.580 -53.940 ;
    END
  END ADC2_OUT[1]
  PIN ADC2_OUT[2]
    PORT
      LAYER met2 ;
        RECT -7.360 -89.860 -7.220 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT -7.450 -63.460 -7.130 -63.140 ;
    END
  END ADC2_OUT[2]
  PIN ADC2_OUT[3]
    PORT
      LAYER met2 ;
        RECT -6.950 -89.860 -6.810 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT -7.010 -81.590 -6.750 -81.270 ;
    END
  END ADC2_OUT[3]
  PIN ADC3_OUT[0]
    PORT
      LAYER met2 ;
        RECT 3.730 -89.780 3.870 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.670 -36.130 3.930 -35.810 ;
    END
  END ADC3_OUT[0]
  PIN ADC3_OUT[1]
    PORT
      LAYER met2 ;
        RECT 4.130 -89.780 4.270 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.070 -54.260 4.330 -53.940 ;
    END
  END ADC3_OUT[1]
  PIN ADC3_OUT[2]
    PORT
      LAYER met2 ;
        RECT 4.550 -89.780 4.690 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.460 -63.460 4.780 -63.140 ;
    END
  END ADC3_OUT[2]
  PIN ADC3_OUT[3]
    PORT
      LAYER met2 ;
        RECT 4.960 -89.780 5.100 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 4.900 -81.590 5.160 -81.270 ;
    END
  END ADC3_OUT[3]
  PIN ADC4_OUT[0]
    PORT
      LAYER met2 ;
        RECT 15.500 -89.950 15.640 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.440 -36.130 15.700 -35.810 ;
    END
  END ADC4_OUT[0]
  PIN ADC4_OUT[1]
    PORT
      LAYER met2 ;
        RECT 15.900 -89.950 16.040 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 15.840 -54.260 16.100 -53.940 ;
    END
  END ADC4_OUT[1]
  PIN ADC4_OUT[2]
    PORT
      LAYER met2 ;
        RECT 16.320 -89.950 16.460 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 16.230 -63.460 16.550 -63.140 ;
    END
  END ADC4_OUT[2]
  PIN ADC4_OUT[3]
    PORT
      LAYER met2 ;
        RECT 16.730 -89.950 16.870 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 16.670 -81.590 16.930 -81.270 ;
    END
  END ADC4_OUT[3]
  PIN ADC5_OUT[0]
    PORT
      LAYER met2 ;
        RECT 27.270 -90.070 27.410 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 27.210 -36.130 27.470 -35.810 ;
    END
  END ADC5_OUT[0]
  PIN ADC5_OUT[1]
    PORT
      LAYER met2 ;
        RECT 27.670 -90.070 27.810 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 27.610 -54.260 27.870 -53.940 ;
    END
  END ADC5_OUT[1]
  PIN ADC5_OUT[2]
    PORT
      LAYER met2 ;
        RECT 28.090 -90.070 28.230 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.000 -63.460 28.320 -63.140 ;
    END
  END ADC5_OUT[2]
  PIN ADC5_OUT[3]
    PORT
      LAYER met2 ;
        RECT 28.500 -90.070 28.640 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.440 -81.590 28.700 -81.270 ;
    END
  END ADC5_OUT[3]
  PIN ADC6_OUT[0]
    PORT
      LAYER met2 ;
        RECT 39.090 -90.180 39.230 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 39.030 -36.130 39.290 -35.810 ;
    END
  END ADC6_OUT[0]
  PIN ADC6_OUT[1]
    PORT
      LAYER met2 ;
        RECT 39.490 -90.180 39.630 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 39.430 -54.260 39.690 -53.940 ;
    END
  END ADC6_OUT[1]
  PIN ADC6_OUT[2]
    PORT
      LAYER met2 ;
        RECT 39.910 -90.180 40.050 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 39.820 -63.460 40.140 -63.140 ;
    END
  END ADC6_OUT[2]
  PIN ADC6_OUT[3]
    PORT
      LAYER met2 ;
        RECT 40.320 -90.180 40.460 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 40.260 -81.590 40.520 -81.270 ;
    END
  END ADC6_OUT[3]
  PIN ADC7_OUT[0]
    PORT
      LAYER met2 ;
        RECT 50.950 -90.260 51.090 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 50.890 -36.130 51.150 -35.810 ;
    END
  END ADC7_OUT[0]
  PIN ADC7_OUT[1]
    PORT
      LAYER met2 ;
        RECT 51.350 -90.260 51.490 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 51.290 -54.260 51.550 -53.940 ;
    END
  END ADC7_OUT[1]
  PIN ADC7_OUT[2]
    PORT
      LAYER met2 ;
        RECT 51.770 -90.260 51.910 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 51.680 -63.460 52.000 -63.140 ;
    END
  END ADC7_OUT[2]
  PIN ADC7_OUT[3]
    PORT
      LAYER met2 ;
        RECT 52.180 -90.260 52.320 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 52.120 -81.590 52.380 -81.270 ;
    END
  END ADC7_OUT[3]
  PIN ADC8_OUT[0]
    PORT
      LAYER met2 ;
        RECT 62.740 -90.230 62.880 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 62.680 -36.130 62.940 -35.810 ;
    END
  END ADC8_OUT[0]
  PIN ADC8_OUT[1]
    PORT
      LAYER met2 ;
        RECT 63.140 -90.230 63.280 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 63.080 -54.260 63.340 -53.940 ;
    END
  END ADC8_OUT[1]
  PIN ADC8_OUT[2]
    PORT
      LAYER met2 ;
        RECT 63.560 -90.230 63.700 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 63.470 -63.460 63.790 -63.140 ;
    END
  END ADC8_OUT[2]
  PIN ADC8_OUT[3]
    PORT
      LAYER met2 ;
        RECT 63.970 -90.230 64.110 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 63.910 -81.590 64.170 -81.270 ;
    END
  END ADC8_OUT[3]
  PIN ADC9_OUT[0]
    PORT
      LAYER met2 ;
        RECT 74.620 -90.120 74.760 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 74.560 -36.130 74.820 -35.810 ;
    END
  END ADC9_OUT[0]
  PIN ADC9_OUT[1]
    PORT
      LAYER met2 ;
        RECT 75.020 -90.120 75.160 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 74.960 -54.260 75.220 -53.940 ;
    END
  END ADC9_OUT[1]
  PIN ADC9_OUT[2]
    PORT
      LAYER met2 ;
        RECT 75.440 -90.120 75.580 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 75.350 -63.460 75.670 -63.140 ;
    END
  END ADC9_OUT[2]
  PIN ADC9_OUT[3]
    PORT
      LAYER met2 ;
        RECT 75.850 -90.120 75.990 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 75.790 -81.590 76.050 -81.270 ;
    END
  END ADC9_OUT[3]
  PIN ADC10_OUT[0]
    PORT
      LAYER met2 ;
        RECT 86.350 -90.270 86.490 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 86.290 -36.130 86.550 -35.810 ;
    END
  END ADC10_OUT[0]
  PIN ADC10_OUT[1]
    PORT
      LAYER met2 ;
        RECT 86.750 -90.270 86.890 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 86.690 -54.260 86.950 -53.940 ;
    END
  END ADC10_OUT[1]
  PIN ADC10_OUT[2]
    PORT
      LAYER met2 ;
        RECT 87.170 -90.270 87.310 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 87.080 -63.460 87.400 -63.140 ;
    END
  END ADC10_OUT[2]
  PIN ADC10_OUT[3]
    PORT
      LAYER met2 ;
        RECT 87.580 -90.270 87.720 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 87.520 -81.590 87.780 -81.270 ;
    END
  END ADC10_OUT[3]
  PIN ADC11_OUT[0]
    PORT
      LAYER met2 ;
        RECT 98.170 -90.350 98.310 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 98.110 -36.130 98.370 -35.810 ;
    END
  END ADC11_OUT[0]
  PIN ADC11_OUT[1]
    PORT
      LAYER met2 ;
        RECT 98.570 -90.350 98.710 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 98.510 -54.260 98.770 -53.940 ;
    END
  END ADC11_OUT[1]
  PIN ADC11_OUT[2]
    PORT
      LAYER met2 ;
        RECT 98.990 -90.350 99.130 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 98.900 -63.460 99.220 -63.140 ;
    END
  END ADC11_OUT[2]
  PIN ADC11_OUT[3]
    PORT
      LAYER met2 ;
        RECT 99.400 -90.350 99.540 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 99.340 -81.590 99.600 -81.270 ;
    END
  END ADC11_OUT[3]
  PIN ADC12_OUT[0]
    PORT
      LAYER met2 ;
        RECT 110.060 -90.170 110.200 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 110.000 -36.130 110.260 -35.810 ;
    END
  END ADC12_OUT[0]
  PIN ADC12_OUT[1]
    PORT
      LAYER met2 ;
        RECT 110.460 -90.170 110.600 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 110.400 -54.260 110.660 -53.940 ;
    END
  END ADC12_OUT[1]
  PIN ADC12_OUT[2]
    PORT
      LAYER met2 ;
        RECT 110.880 -90.170 111.020 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 110.790 -63.460 111.110 -63.140 ;
    END
  END ADC12_OUT[2]
  PIN ADC12_OUT[3]
    PORT
      LAYER met2 ;
        RECT 111.290 -90.170 111.430 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 111.230 -81.590 111.490 -81.270 ;
    END
  END ADC12_OUT[3]
  PIN ADC13_OUT[0]
    PORT
      LAYER met2 ;
        RECT 122.010 -90.130 122.150 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 121.950 -36.130 122.210 -35.810 ;
    END
  END ADC13_OUT[0]
  PIN ADC13_OUT[1]
    PORT
      LAYER met2 ;
        RECT 122.410 -90.130 122.550 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 122.350 -54.260 122.610 -53.940 ;
    END
  END ADC13_OUT[1]
  PIN ADC13_OUT[2]
    PORT
      LAYER met2 ;
        RECT 122.830 -90.130 122.970 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 122.740 -63.460 123.060 -63.140 ;
    END
  END ADC13_OUT[2]
  PIN ADC13_OUT[3]
    PORT
      LAYER met2 ;
        RECT 123.240 -90.130 123.380 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 123.180 -81.590 123.440 -81.270 ;
    END
  END ADC13_OUT[3]
  PIN ADC14_OUT[0]
    PORT
      LAYER met2 ;
        RECT 133.770 -90.070 133.910 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 133.710 -36.130 133.970 -35.810 ;
    END
  END ADC14_OUT[0]
  PIN ADC14_OUT[1]
    PORT
      LAYER met2 ;
        RECT 134.170 -90.070 134.310 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 134.110 -54.260 134.370 -53.940 ;
    END
  END ADC14_OUT[1]
  PIN ADC14_OUT[2]
    PORT
      LAYER met2 ;
        RECT 134.590 -90.070 134.730 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 134.500 -63.460 134.820 -63.140 ;
    END
  END ADC14_OUT[2]
  PIN ADC14_OUT[3]
    PORT
      LAYER met2 ;
        RECT 135.000 -90.070 135.140 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 134.940 -81.590 135.200 -81.270 ;
    END
  END ADC14_OUT[3]
  PIN ADC15_OUT[0]
    PORT
      LAYER met2 ;
        RECT 142.810 -90.110 142.950 -36.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 142.750 -36.130 143.010 -35.810 ;
    END
  END ADC15_OUT[0]
  PIN ADC15_OUT[1]
    PORT
      LAYER met2 ;
        RECT 143.210 -90.110 143.350 -54.260 ;
    END
    PORT
      LAYER met2 ;
        RECT 143.150 -54.260 143.410 -53.940 ;
    END
  END ADC15_OUT[1]
  PIN ADC15_OUT[2]
    PORT
      LAYER met2 ;
        RECT 143.630 -90.110 143.770 -63.460 ;
    END
    PORT
      LAYER met2 ;
        RECT 143.540 -63.460 143.860 -63.140 ;
    END
  END ADC15_OUT[2]
  PIN ADC15_OUT[3]
    PORT
      LAYER met2 ;
        RECT 144.040 -90.110 144.180 -81.590 ;
    END
    PORT
      LAYER met2 ;
        RECT 143.980 -81.590 144.240 -81.270 ;
    END
  END ADC15_OUT[3]
  PIN Din[0]
    PORT
      LAYER met2 ;
        RECT 2.250 -21.300 2.570 -20.980 ;
    END
    PORT
      LAYER met2 ;
        RECT 2.340 -20.980 2.480 53.560 ;
    END
  END Din[0]
  PIN Din[1]
    PORT
      LAYER met2 ;
        RECT 8.060 -21.280 8.380 -20.960 ;
    END
    PORT
      LAYER met2 ;
        RECT 8.150 -20.960 8.290 53.450 ;
    END
  END Din[1]
  PIN Din[2]
    PORT
      LAYER met2 ;
        RECT 13.780 -21.290 14.100 -20.970 ;
    END
    PORT
      LAYER met2 ;
        RECT 13.860 -20.970 14.000 53.410 ;
    END
  END Din[2]
  PIN Din[3]
    PORT
      LAYER met2 ;
        RECT 19.560 -21.310 19.880 -20.990 ;
    END
    PORT
      LAYER met2 ;
        RECT 19.640 -20.990 19.780 53.420 ;
    END
  END Din[3]
  PIN Din[4]
    PORT
      LAYER met2 ;
        RECT 25.310 -21.310 25.630 -20.990 ;
    END
    PORT
      LAYER met2 ;
        RECT 25.370 -20.990 25.510 53.420 ;
    END
  END Din[4]
  PIN Din[5]
    PORT
      LAYER met2 ;
        RECT 31.020 -21.330 31.340 -21.010 ;
    END
    PORT
      LAYER met2 ;
        RECT 31.100 -21.010 31.240 53.400 ;
    END
  END Din[5]
  PIN Din[6]
    PORT
      LAYER met2 ;
        RECT 36.790 -21.320 37.110 -21.000 ;
    END
    PORT
      LAYER met2 ;
        RECT 36.860 -21.000 37.000 53.410 ;
    END
  END Din[6]
  PIN Din[7]
    PORT
      LAYER met2 ;
        RECT 42.590 -21.310 42.910 -20.990 ;
    END
    PORT
      LAYER met2 ;
        RECT 42.640 -20.990 42.780 53.420 ;
    END
  END Din[7]
  PIN Din[8]
    PORT
      LAYER met2 ;
        RECT 48.290 -21.300 48.610 -20.980 ;
    END
    PORT
      LAYER met2 ;
        RECT 48.370 -20.980 48.510 53.420 ;
    END
  END Din[8]
  PIN Din[9]
    PORT
      LAYER met2 ;
        RECT 54.060 -21.320 54.380 -21.000 ;
    END
    PORT
      LAYER met2 ;
        RECT 54.120 -21.000 54.260 53.400 ;
    END
  END Din[9]
  PIN Din[10]
    PORT
      LAYER met2 ;
        RECT 59.800 -21.300 60.120 -20.980 ;
    END
    PORT
      LAYER met2 ;
        RECT 59.880 -20.980 60.020 53.410 ;
    END
  END Din[10]
  PIN Din[11]
    PORT
      LAYER met2 ;
        RECT 65.530 -21.310 65.850 -20.990 ;
    END
    PORT
      LAYER met2 ;
        RECT 65.610 -20.990 65.750 53.410 ;
    END
  END Din[11]
  PIN Din[12]
    PORT
      LAYER met2 ;
        RECT 71.300 -21.320 71.620 -21.000 ;
    END
    PORT
      LAYER met2 ;
        RECT 71.360 -21.000 71.500 53.410 ;
    END
  END Din[12]
  PIN Din[13]
    PORT
      LAYER met2 ;
        RECT 77.060 -21.320 77.380 -21.000 ;
    END
    PORT
      LAYER met2 ;
        RECT 77.110 -21.000 77.250 53.420 ;
    END
  END Din[13]
  PIN Din[14]
    PORT
      LAYER met2 ;
        RECT 82.790 -21.340 83.110 -21.020 ;
    END
    PORT
      LAYER met2 ;
        RECT 82.880 -21.020 83.020 53.420 ;
    END
  END Din[14]
  PIN Din[15]
    PORT
      LAYER met2 ;
        RECT 88.540 -21.340 88.860 -21.020 ;
    END
    PORT
      LAYER met2 ;
        RECT 88.630 -21.020 88.770 53.420 ;
    END
  END Din[15]
  PIN WWLD[0]
    PORT
      LAYER met1 ;
        RECT 92.300 47.090 92.590 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 47.090 86.840 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 47.090 81.090 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 47.090 75.340 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 47.090 69.590 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 47.090 63.840 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 47.090 58.090 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 47.090 52.340 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 47.090 46.590 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 47.090 40.840 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 47.090 35.090 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 47.090 29.340 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 47.090 23.590 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 47.090 17.840 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 47.090 12.090 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 47.090 6.340 47.210 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 47.210 94.660 47.350 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 47.350 90.980 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 47.350 85.230 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 47.350 79.480 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 47.350 73.730 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 47.350 67.980 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 47.350 62.230 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 47.350 56.480 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 47.350 50.730 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 47.350 44.980 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 47.350 39.230 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 47.350 33.480 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 47.350 27.730 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 47.350 21.980 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 47.350 16.230 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 47.350 10.480 47.470 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 47.350 4.730 47.470 ;
    END
  END WWLD[0]
  PIN WWLD[1]
    PORT
      LAYER met1 ;
        RECT 92.300 44.680 92.590 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 44.680 86.840 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 44.680 81.090 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 44.680 75.340 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 44.680 69.590 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 44.680 63.840 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 44.680 58.090 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 44.680 52.340 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 44.680 46.590 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 44.680 40.840 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 44.680 35.090 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 44.680 29.340 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 44.680 23.590 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 44.680 17.840 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 44.680 12.090 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 44.680 6.340 44.800 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 44.800 94.660 44.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 44.940 90.980 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 44.940 85.230 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 44.940 79.480 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 44.940 73.730 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 44.940 67.980 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 44.940 62.230 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 44.940 56.480 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 44.940 50.730 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 44.940 44.980 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 44.940 39.230 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 44.940 33.480 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 44.940 27.730 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 44.940 21.980 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 44.940 16.230 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 44.940 10.480 45.060 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 44.940 4.730 45.060 ;
    END
  END WWLD[1]
  PIN WWLD[2]
    PORT
      LAYER met1 ;
        RECT 92.300 41.710 92.590 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 41.710 86.840 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 41.710 81.090 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 41.710 75.340 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 41.710 69.590 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 41.710 63.840 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 41.710 58.090 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 41.710 52.340 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 41.710 46.590 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 41.710 40.840 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 41.710 35.090 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 41.710 29.340 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 41.710 23.590 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 41.710 17.840 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 41.710 12.090 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 41.710 6.340 41.830 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 41.830 94.660 41.970 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 41.970 90.980 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 41.970 85.230 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 41.970 79.480 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 41.970 73.730 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 41.970 67.980 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 41.970 62.230 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 41.970 56.480 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 41.970 50.730 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 41.970 44.980 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 41.970 39.230 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 41.970 33.480 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 41.970 27.730 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 41.970 21.980 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 41.970 16.230 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 41.970 10.480 42.090 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 41.970 4.730 42.090 ;
    END
  END WWLD[2]
  PIN WWLD[3]
    PORT
      LAYER met1 ;
        RECT 92.300 39.300 92.590 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 39.300 86.840 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 39.300 81.090 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 39.300 75.340 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 39.300 69.590 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 39.300 63.840 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 39.300 58.090 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 39.300 52.340 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 39.300 46.590 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 39.300 40.840 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 39.300 35.090 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 39.300 29.340 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 39.300 23.590 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 39.300 17.840 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 39.300 12.090 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 39.300 6.340 39.420 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 39.420 94.660 39.560 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 39.560 90.980 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 39.560 85.230 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 39.560 79.480 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 39.560 73.730 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 39.560 67.980 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 39.560 62.230 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 39.560 56.480 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 39.560 50.730 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 39.560 44.980 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 39.560 39.230 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 39.560 33.480 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 39.560 27.730 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 39.560 21.980 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 39.560 16.230 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 39.560 10.480 39.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 39.560 4.730 39.680 ;
    END
  END WWLD[3]
  PIN WWLD[4]
    PORT
      LAYER met1 ;
        RECT 92.300 -2.480 92.590 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 -2.480 86.840 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 -2.480 81.090 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 -2.480 75.340 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 -2.480 69.590 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 -2.480 63.840 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 -2.480 58.090 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 -2.480 52.340 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 -2.480 46.590 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 -2.480 40.840 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 -2.480 35.090 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 -2.480 29.340 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 -2.480 23.590 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 -2.480 17.840 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 -2.480 12.090 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 -2.480 6.340 -2.360 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 -2.360 94.660 -2.220 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 -2.220 90.980 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 -2.220 85.230 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 -2.220 79.480 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 -2.220 73.730 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 -2.220 67.980 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 -2.220 62.230 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 -2.220 56.480 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 -2.220 50.730 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 -2.220 44.980 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 -2.220 39.230 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 -2.220 33.480 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 -2.220 27.730 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 -2.220 21.980 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 -2.220 16.230 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 -2.220 10.480 -2.100 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 -2.220 4.730 -2.100 ;
    END
  END WWLD[4]
  PIN WWLD[5]
    PORT
      LAYER met1 ;
        RECT 92.300 -4.890 92.590 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 -4.890 86.840 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 -4.890 81.090 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 -4.890 75.340 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 -4.890 69.590 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 -4.890 63.840 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 -4.890 58.090 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 -4.890 52.340 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 -4.890 46.590 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 -4.890 40.840 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 -4.890 35.090 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 -4.890 29.340 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 -4.890 23.590 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 -4.890 17.840 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 -4.890 12.090 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 -4.890 6.340 -4.770 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 -4.770 94.660 -4.630 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 -4.630 90.980 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 -4.630 85.230 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 -4.630 79.480 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 -4.630 73.730 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 -4.630 67.980 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 -4.630 62.230 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 -4.630 56.480 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 -4.630 50.730 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 -4.630 44.980 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 -4.630 39.230 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 -4.630 33.480 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 -4.630 27.730 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 -4.630 21.980 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 -4.630 16.230 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 -4.630 10.480 -4.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 -4.630 4.730 -4.510 ;
    END
  END WWLD[5]
  PIN WWLD[6]
    PORT
      LAYER met1 ;
        RECT 92.300 -7.890 92.590 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 -7.890 86.840 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 -7.890 81.090 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 -7.890 75.340 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 -7.890 69.590 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 -7.890 63.840 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 -7.890 58.090 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 -7.890 52.340 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 -7.890 46.590 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 -7.890 40.840 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 -7.890 35.090 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 -7.890 29.340 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 -7.890 23.590 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 -7.890 17.840 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 -7.890 12.090 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 -7.890 6.340 -7.770 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 -7.770 94.660 -7.630 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 -7.630 90.980 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 -7.630 85.230 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 -7.630 79.480 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 -7.630 73.730 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 -7.630 67.980 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 -7.630 62.230 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 -7.630 56.480 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 -7.630 50.730 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 -7.630 44.980 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 -7.630 39.230 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 -7.630 33.480 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 -7.630 27.730 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 -7.630 21.980 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 -7.630 16.230 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 -7.630 10.480 -7.510 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 -7.630 4.730 -7.510 ;
    END
  END WWLD[6]
  PIN WWLD[7]
    PORT
      LAYER met1 ;
        RECT 92.300 -10.300 92.590 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 86.550 -10.300 86.840 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 80.800 -10.300 81.090 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 75.050 -10.300 75.340 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.300 -10.300 69.590 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 63.550 -10.300 63.840 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 57.800 -10.300 58.090 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 52.050 -10.300 52.340 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 46.300 -10.300 46.590 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 40.550 -10.300 40.840 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 34.800 -10.300 35.090 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 29.050 -10.300 29.340 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 23.300 -10.300 23.590 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.550 -10.300 17.840 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.800 -10.300 12.090 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.050 -10.300 6.340 -10.180 ;
    END
    PORT
      LAYER met1 ;
        RECT -45.490 -10.180 94.660 -10.040 ;
    END
    PORT
      LAYER met1 ;
        RECT 90.690 -10.040 90.980 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 84.940 -10.040 85.230 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.190 -10.040 79.480 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 73.440 -10.040 73.730 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 67.690 -10.040 67.980 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 61.940 -10.040 62.230 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 56.190 -10.040 56.480 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 50.440 -10.040 50.730 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 44.690 -10.040 44.980 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.940 -10.040 39.230 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 33.190 -10.040 33.480 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.440 -10.040 27.730 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 21.690 -10.040 21.980 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 15.940 -10.040 16.230 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 10.190 -10.040 10.480 -9.920 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.440 -10.040 4.730 -9.920 ;
    END
  END WWLD[7]
  PIN SA_OUT[0]
    PORT
      LAYER met3 ;
        RECT 5.930 -6.400 6.290 -6.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.930 -6.370 100.480 -6.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.930 -6.070 6.290 -6.040 ;
    END
  END SA_OUT[0]
  PIN SA_OUT[1]
    PORT
      LAYER met3 ;
        RECT 11.680 -7.670 12.040 -7.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.680 -7.640 100.480 -7.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.680 -7.340 12.040 -7.310 ;
    END
  END SA_OUT[1]
  PIN SA_OUT[2]
    PORT
      LAYER met3 ;
        RECT 17.480 -9.040 17.840 -9.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.480 -9.010 100.480 -8.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.480 -8.710 17.840 -8.680 ;
    END
  END SA_OUT[2]
  PIN SA_OUT[3]
    PORT
      LAYER met3 ;
        RECT 23.180 -10.210 23.540 -10.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.180 -10.180 100.480 -9.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.180 -9.880 23.540 -9.850 ;
    END
  END SA_OUT[3]
  PIN SA_OUT[4]
    PORT
      LAYER met3 ;
        RECT 28.930 -11.460 29.290 -11.430 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.930 -11.430 100.480 -11.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.930 -11.130 29.290 -11.100 ;
    END
  END SA_OUT[4]
  PIN SA_OUT[5]
    PORT
      LAYER met3 ;
        RECT 34.680 -12.910 35.040 -12.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.680 -12.880 100.480 -12.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.680 -12.580 35.040 -12.550 ;
    END
  END SA_OUT[5]
  PIN SA_OUT[6]
    PORT
      LAYER met3 ;
        RECT 40.400 -14.150 40.800 -14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.400 -14.100 100.480 -13.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.400 -13.800 40.800 -13.750 ;
    END
  END SA_OUT[6]
  PIN SA_OUT[7]
    PORT
      LAYER met3 ;
        RECT 46.180 -15.010 46.540 -14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.180 -14.980 100.480 -14.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.180 -14.680 46.540 -14.650 ;
    END
  END SA_OUT[7]
  PIN SA_OUT[8]
    PORT
      LAYER met3 ;
        RECT 51.930 -15.840 52.290 -15.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.930 -15.810 100.480 -15.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.930 -15.510 52.290 -15.480 ;
    END
  END SA_OUT[8]
  PIN SA_OUT[9]
    PORT
      LAYER met3 ;
        RECT 57.680 -16.620 58.040 -16.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.680 -16.590 100.480 -16.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.680 -16.290 58.040 -16.260 ;
    END
  END SA_OUT[9]
  PIN SA_OUT[10]
    PORT
      LAYER met3 ;
        RECT 63.430 -17.480 63.790 -17.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 -17.450 100.480 -17.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 -17.150 63.790 -17.120 ;
    END
  END SA_OUT[10]
  PIN SA_OUT[11]
    PORT
      LAYER met3 ;
        RECT 69.180 -18.280 69.540 -18.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.180 -18.250 100.480 -17.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.180 -17.950 69.540 -17.920 ;
    END
  END SA_OUT[11]
  PIN SA_OUT[12]
    PORT
      LAYER met3 ;
        RECT 74.930 -19.080 75.290 -19.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.930 -19.050 100.480 -18.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.930 -18.750 75.290 -18.720 ;
    END
  END SA_OUT[12]
  PIN SA_OUT[13]
    PORT
      LAYER met3 ;
        RECT 80.680 -19.730 81.040 -19.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.680 -19.700 100.480 -19.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.680 -19.400 81.040 -19.370 ;
    END
  END SA_OUT[13]
  PIN SA_OUT[14]
    PORT
      LAYER met3 ;
        RECT 86.430 -20.870 86.790 -20.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.430 -20.840 100.480 -20.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.430 -20.540 86.790 -20.510 ;
    END
  END SA_OUT[14]
  PIN SA_OUT[15]
    PORT
      LAYER met3 ;
        RECT 92.180 -21.760 92.540 -21.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.180 -21.730 100.480 -21.430 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.180 -21.430 92.540 -21.400 ;
    END
  END SA_OUT[15]
  PIN EN
    PORT
      LAYER met3 ;
        RECT 89.320 -24.540 89.720 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.800 -24.540 88.200 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.840 -24.540 78.240 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.310 -24.540 76.710 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 -24.550 66.730 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.800 -24.550 65.200 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.840 -24.540 55.240 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.290 -24.540 53.690 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.360 -24.550 43.760 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.770 -24.540 42.170 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.840 -24.540 32.240 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.300 -24.540 30.700 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.350 -24.540 20.750 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.800 -24.540 19.200 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.850 -24.540 9.250 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.300 -24.540 7.700 -24.490 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.420 -24.490 89.720 -24.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.320 -24.190 89.720 -24.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.800 -24.190 88.200 -24.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.840 -24.190 78.240 -24.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.310 -24.190 76.710 -24.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 -24.190 66.730 -24.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.800 -24.190 65.200 -24.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.840 -24.190 55.240 -24.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.290 -24.190 53.690 -24.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.360 -24.190 43.760 -24.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.770 -24.190 42.170 -24.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.840 -24.190 32.240 -24.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.300 -24.190 30.700 -24.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.350 -24.190 20.750 -24.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.800 -24.190 19.200 -24.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.850 -24.190 9.250 -24.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.300 -24.190 7.700 -24.140 ;
    END
  END EN
  PIN PRE_A
    PORT
      LAYER met3 ;
        RECT 85.110 -25.290 85.510 -25.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.530 -25.300 80.930 -25.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.610 -25.270 74.010 -25.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.030 -25.270 69.430 -25.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.540 -25.270 57.940 -25.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.030 -25.310 46.430 -25.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.120 -25.290 39.520 -25.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.540 -25.270 34.940 -25.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.620 -25.290 28.020 -25.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.030 -25.280 23.430 -25.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 -25.310 5.010 -25.250 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.420 -25.250 92.390 -24.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.030 -24.950 92.390 -24.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.110 -24.950 85.510 -24.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.530 -24.950 80.930 -24.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.610 -24.950 74.010 -24.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.030 -24.950 69.430 -24.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.110 -24.950 62.510 -24.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.540 -24.950 57.940 -24.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.610 -24.950 51.010 -24.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.030 -24.950 46.430 -24.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.120 -24.950 39.520 -24.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.540 -24.950 34.940 -24.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.620 -24.950 28.020 -24.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.030 -24.950 23.430 -24.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.100 -24.950 16.500 -24.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.540 -24.950 11.940 -24.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 -24.950 5.010 -24.910 ;
    END
  END PRE_A
  PIN VDD
    PORT
      LAYER met3 ;
        RECT 139.020 -31.030 139.380 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.010 -31.010 130.370 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.140 -30.990 118.500 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.270 -31.030 106.630 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.430 -31.020 94.790 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.590 -31.010 82.950 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.770 -31.030 71.130 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.950 -31.030 59.310 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.130 -31.000 47.490 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.310 -31.030 35.670 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.490 -31.030 23.850 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.670 -31.020 12.030 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.140 -31.040 0.220 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.770 -31.000 -23.410 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.270 -31.000 -34.910 -30.970 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.150 -30.970 144.360 -30.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.010 -30.670 130.370 -30.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.140 -30.670 118.500 -30.630 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.430 -30.670 94.790 -30.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.590 -30.670 82.950 -30.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.130 -30.670 47.490 -30.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.670 -30.670 12.030 -30.660 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.770 -30.670 -23.410 -30.640 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.270 -30.670 -34.910 -30.640 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.170 -30.670 -42.810 -30.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.690 50.330 63.090 50.340 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.170 50.280 -42.810 50.340 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.490 50.340 100.380 50.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.420 50.640 91.820 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.670 50.640 86.070 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.930 50.640 80.330 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.180 50.640 74.580 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.430 50.640 68.830 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.690 50.640 63.090 50.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.940 50.640 57.340 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.180 50.640 51.580 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.430 50.640 45.830 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.680 50.640 40.080 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.930 50.640 34.330 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.190 50.640 28.590 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 50.640 22.830 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.700 50.640 17.100 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 50.640 11.350 50.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.190 50.640 5.590 50.740 ;
    END
    PORT
      LAYER nwell ;
        RECT 135.850 -86.240 142.470 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 126.840 -86.240 133.460 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 114.970 -86.240 121.590 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 103.100 -86.240 109.720 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 91.260 -86.240 97.880 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 79.420 -86.240 86.040 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 67.600 -86.240 74.220 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 55.780 -86.240 62.400 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 43.960 -86.240 50.580 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 32.140 -86.240 38.760 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 20.320 -86.240 26.940 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 8.500 -86.240 15.120 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT -3.310 -86.240 3.310 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT -26.940 -86.240 -20.320 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT -38.440 -86.240 -31.820 -81.270 ;
    END
    PORT
      LAYER nwell ;
        RECT 135.850 -63.470 142.470 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 126.840 -63.470 133.460 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 114.970 -63.470 121.590 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 103.100 -63.470 109.720 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 91.260 -63.470 97.880 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 79.420 -63.470 86.040 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 67.600 -63.470 74.220 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 55.780 -63.470 62.400 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 43.960 -63.470 50.580 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 32.140 -63.470 38.760 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 20.320 -63.470 26.940 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 8.500 -63.470 15.120 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT -3.310 -63.470 3.310 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT -26.940 -63.470 -20.320 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT -38.440 -63.470 -31.820 -53.940 ;
    END
    PORT
      LAYER nwell ;
        RECT 135.850 -36.140 142.470 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 126.840 -36.140 133.460 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 114.970 -36.140 121.590 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 103.100 -36.140 109.720 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 91.260 -36.140 97.880 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 79.420 -36.140 86.040 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 67.600 -36.140 74.220 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 55.780 -36.140 62.400 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 43.960 -36.140 50.580 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 32.140 -36.140 38.760 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 20.320 -36.140 26.940 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 8.500 -36.140 15.120 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT -3.310 -36.140 3.310 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT -26.940 -36.140 -20.320 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT -38.440 -36.140 -31.820 -31.170 ;
    END
    PORT
      LAYER nwell ;
        RECT 91.140 -24.540 94.660 -21.210 ;
    END
    PORT
      LAYER nwell ;
        RECT 79.640 -24.540 86.390 -21.210 ;
    END
    PORT
      LAYER nwell ;
        RECT 68.140 -24.540 74.890 -21.210 ;
    END
    PORT
      LAYER nwell ;
        RECT 56.640 -24.540 63.390 -21.210 ;
    END
    PORT
      LAYER nwell ;
        RECT 45.140 -24.540 51.890 -21.210 ;
    END
    PORT
      LAYER nwell ;
        RECT 33.640 -24.540 40.390 -21.210 ;
    END
    PORT
      LAYER nwell ;
        RECT 22.140 -24.540 28.890 -21.210 ;
    END
    PORT
      LAYER nwell ;
        RECT 10.640 -24.540 17.390 -21.210 ;
    END
    PORT
      LAYER nwell ;
        RECT 2.250 -24.540 5.890 -21.210 ;
    END
    PORT
      LAYER nwell ;
        RECT 2.250 -14.140 94.660 -11.420 ;
    END
    PORT
      LAYER nwell ;
        RECT 90.950 -11.420 92.330 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 85.200 -11.420 86.580 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 79.450 -11.420 80.830 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 73.700 -11.420 75.080 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 67.950 -11.420 69.330 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 62.200 -11.420 63.580 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 56.450 -11.420 57.830 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 50.700 -11.420 52.080 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 44.950 -11.420 46.330 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 39.200 -11.420 40.580 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 33.450 -11.420 34.830 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 27.700 -11.420 29.080 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 21.950 -11.420 23.330 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 16.200 -11.420 17.580 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 10.450 -11.420 11.830 50.590 ;
    END
    PORT
      LAYER nwell ;
        RECT 4.700 -11.420 6.080 50.590 ;
    END
  END VDD
  PIN VSS
    PORT
      LAYER met3 ;
        RECT 88.650 -23.540 89.050 -23.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.080 -23.560 77.480 -23.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.630 -23.560 66.030 -23.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.950 -23.560 54.350 -23.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.550 -23.580 42.950 -23.530 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.540 -23.530 42.950 -23.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.980 -23.570 31.380 -23.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.970 -23.520 31.380 -23.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.550 -23.560 19.950 -23.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.060 -23.550 8.460 -23.510 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.350 -23.510 89.050 -23.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.640 -23.210 89.050 -23.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.650 -23.190 89.050 -23.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.080 -23.210 77.480 -23.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.630 -23.210 66.030 -23.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.950 -23.210 54.350 -23.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.550 -23.210 42.950 -23.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.980 -23.210 31.380 -23.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.550 -23.210 19.950 -23.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.050 -23.210 8.460 -23.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.060 -23.200 8.460 -23.150 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.350 -23.210 -0.050 -20.650 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.400 -20.650 0.000 -20.600 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.830 -20.670 -41.470 -20.600 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.520 -20.600 0.000 -20.300 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.400 -20.300 0.000 -20.250 ;
    END
    PORT
      LAYER pwell ;
        RECT 135.850 -81.270 142.470 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 126.840 -81.270 133.460 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 114.970 -81.270 121.590 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 103.100 -81.270 109.720 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 91.260 -81.270 97.880 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 79.420 -81.270 86.040 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 67.600 -81.270 74.220 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 55.780 -81.270 62.400 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 43.960 -81.270 50.580 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 32.140 -81.270 38.760 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 20.320 -81.270 26.940 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 8.500 -81.270 15.120 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT -3.310 -81.270 3.310 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT -15.120 -81.270 -8.500 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT -26.940 -81.270 -20.320 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT -38.440 -81.270 -31.820 -63.470 ;
    END
    PORT
      LAYER pwell ;
        RECT 135.850 -53.940 142.470 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 126.840 -53.940 133.460 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 114.970 -53.940 121.590 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 103.100 -53.940 109.720 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 91.260 -53.940 97.880 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 79.420 -53.940 86.040 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 67.600 -53.940 74.220 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 55.780 -53.940 62.400 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 43.960 -53.940 50.580 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 32.140 -53.940 38.760 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 20.320 -53.940 26.940 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 8.500 -53.940 15.120 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT -3.310 -53.940 3.310 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT -15.120 -53.940 -8.500 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT -26.940 -53.940 -20.320 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT -38.440 -53.940 -31.820 -36.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 86.390 -24.540 91.140 -22.560 ;
    END
    PORT
      LAYER pwell ;
        RECT 74.890 -24.540 79.640 -22.560 ;
    END
    PORT
      LAYER pwell ;
        RECT 63.390 -24.540 68.140 -22.560 ;
    END
    PORT
      LAYER pwell ;
        RECT 51.890 -24.540 56.640 -22.560 ;
    END
    PORT
      LAYER pwell ;
        RECT 40.390 -24.540 45.140 -22.560 ;
    END
    PORT
      LAYER pwell ;
        RECT 28.890 -24.540 33.640 -22.560 ;
    END
    PORT
      LAYER pwell ;
        RECT 17.390 -24.540 22.140 -22.560 ;
    END
    PORT
      LAYER pwell ;
        RECT 5.890 -24.540 10.640 -22.560 ;
    END
    PORT
      LAYER pwell ;
        RECT 2.250 -21.210 94.660 -14.140 ;
    END
    PORT
      LAYER pwell ;
        RECT 92.330 -11.420 94.660 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 86.580 -11.420 90.950 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 80.830 -11.420 85.200 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 75.080 -11.420 79.450 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 69.330 -11.420 73.700 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 63.580 -11.420 67.950 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 57.830 -11.420 62.200 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 52.080 -11.420 56.450 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 46.330 -11.420 50.700 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 40.580 -11.420 44.950 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 34.830 -11.420 39.200 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 29.080 -11.420 33.450 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 23.330 -11.420 27.700 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 17.580 -11.420 21.950 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 11.830 -11.420 16.200 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 6.080 -11.420 10.450 48.670 ;
    END
    PORT
      LAYER pwell ;
        RECT 2.250 -11.420 4.700 48.670 ;
    END
  END VSS
  PIN Iref0
    PORT
      LAYER met2 ;
        RECT 144.510 -90.100 144.680 -44.740 ;
    END
    PORT
      LAYER met2 ;
        RECT 144.460 -44.740 144.720 -44.420 ;
    END
  END Iref0
  PIN Iref1
    PORT
      LAYER met2 ;
        RECT 145.070 -90.100 145.240 -45.630 ;
    END
    PORT
      LAYER met2 ;
        RECT 145.020 -45.630 145.280 -45.310 ;
    END
  END Iref1
  PIN Iref2
    PORT
      LAYER met2 ;
        RECT 145.610 -90.100 145.780 -72.000 ;
    END
    PORT
      LAYER met2 ;
        RECT 145.560 -72.000 145.820 -71.680 ;
    END
  END Iref2
  PIN Iref3
    PORT
      LAYER met2 ;
        RECT 146.160 -90.100 146.330 -72.970 ;
    END
    PORT
      LAYER met2 ;
        RECT 146.110 -72.970 146.370 -72.650 ;
    END
  END Iref3
  OBS
      LAYER li1 ;
        RECT -43.520 -23.510 146.400 50.950 ;
      LAYER li1 ;
        RECT -43.520 -87.220 147.150 -23.510 ;
      LAYER met1 ;
        RECT -45.490 50.470 146.400 50.950 ;
        RECT -45.490 50.420 4.060 50.470 ;
        RECT 6.690 50.420 9.810 50.470 ;
        RECT 12.440 50.420 15.560 50.470 ;
        RECT 18.190 50.420 21.310 50.470 ;
        RECT 23.940 50.420 27.060 50.470 ;
        RECT 29.690 50.420 32.810 50.470 ;
        RECT 35.440 50.420 38.560 50.470 ;
        RECT 41.190 50.420 44.310 50.470 ;
        RECT 46.940 50.420 50.060 50.470 ;
        RECT 52.690 50.420 55.810 50.470 ;
        RECT 58.440 50.420 61.560 50.470 ;
        RECT 64.190 50.420 67.310 50.470 ;
        RECT 69.940 50.420 73.060 50.470 ;
        RECT 75.690 50.420 78.810 50.470 ;
        RECT 81.440 50.420 84.560 50.470 ;
        RECT 87.190 50.420 90.310 50.470 ;
        RECT 92.940 50.420 146.400 50.470 ;
        RECT 94.940 49.720 146.400 50.420 ;
        RECT -45.490 49.680 4.060 49.720 ;
        RECT 6.690 49.680 9.810 49.720 ;
        RECT 12.440 49.680 15.560 49.720 ;
        RECT 18.190 49.680 21.310 49.720 ;
        RECT 23.940 49.680 27.060 49.720 ;
        RECT 29.690 49.680 32.810 49.720 ;
        RECT 35.440 49.680 38.560 49.720 ;
        RECT 41.190 49.680 44.310 49.720 ;
        RECT 46.940 49.680 50.060 49.720 ;
        RECT 52.690 49.680 55.810 49.720 ;
        RECT 58.440 49.680 61.560 49.720 ;
        RECT 64.190 49.680 67.310 49.720 ;
        RECT 69.940 49.680 73.060 49.720 ;
        RECT 75.690 49.680 78.810 49.720 ;
        RECT 81.440 49.680 84.560 49.720 ;
        RECT 87.190 49.680 90.310 49.720 ;
        RECT 92.940 49.680 146.400 49.720 ;
        RECT -45.490 47.750 146.400 49.680 ;
        RECT -45.490 47.630 4.160 47.750 ;
        RECT 5.010 47.630 9.910 47.750 ;
        RECT 10.760 47.630 15.660 47.750 ;
        RECT 16.510 47.630 21.410 47.750 ;
        RECT 22.260 47.630 27.160 47.750 ;
        RECT 28.010 47.630 32.910 47.750 ;
        RECT 33.760 47.630 38.660 47.750 ;
        RECT 39.510 47.630 44.410 47.750 ;
        RECT 45.260 47.630 50.160 47.750 ;
        RECT 51.010 47.630 55.910 47.750 ;
        RECT 56.760 47.630 61.660 47.750 ;
        RECT 62.510 47.630 67.410 47.750 ;
        RECT 68.260 47.630 73.160 47.750 ;
        RECT 74.010 47.630 78.910 47.750 ;
        RECT 79.760 47.630 84.660 47.750 ;
        RECT 85.510 47.630 90.410 47.750 ;
        RECT 91.260 47.630 146.400 47.750 ;
        RECT 94.940 46.930 146.400 47.630 ;
        RECT -45.490 46.810 5.770 46.930 ;
        RECT 6.620 46.810 11.520 46.930 ;
        RECT 12.370 46.810 17.270 46.930 ;
        RECT 18.120 46.810 23.020 46.930 ;
        RECT 23.870 46.810 28.770 46.930 ;
        RECT 29.620 46.810 34.520 46.930 ;
        RECT 35.370 46.810 40.270 46.930 ;
        RECT 41.120 46.810 46.020 46.930 ;
        RECT 46.870 46.810 51.770 46.930 ;
        RECT 52.620 46.810 57.520 46.930 ;
        RECT 58.370 46.810 63.270 46.930 ;
        RECT 64.120 46.810 69.020 46.930 ;
        RECT 69.870 46.810 74.770 46.930 ;
        RECT 75.620 46.810 80.520 46.930 ;
        RECT 81.370 46.810 86.270 46.930 ;
        RECT 87.120 46.810 92.020 46.930 ;
        RECT 92.870 46.810 146.400 46.930 ;
        RECT -45.490 45.340 146.400 46.810 ;
        RECT -45.490 45.220 4.160 45.340 ;
        RECT 5.010 45.220 9.910 45.340 ;
        RECT 10.760 45.220 15.660 45.340 ;
        RECT 16.510 45.220 21.410 45.340 ;
        RECT 22.260 45.220 27.160 45.340 ;
        RECT 28.010 45.220 32.910 45.340 ;
        RECT 33.760 45.220 38.660 45.340 ;
        RECT 39.510 45.220 44.410 45.340 ;
        RECT 45.260 45.220 50.160 45.340 ;
        RECT 51.010 45.220 55.910 45.340 ;
        RECT 56.760 45.220 61.660 45.340 ;
        RECT 62.510 45.220 67.410 45.340 ;
        RECT 68.260 45.220 73.160 45.340 ;
        RECT 74.010 45.220 78.910 45.340 ;
        RECT 79.760 45.220 84.660 45.340 ;
        RECT 85.510 45.220 90.410 45.340 ;
        RECT 91.260 45.220 146.400 45.340 ;
        RECT 94.940 44.520 146.400 45.220 ;
        RECT -45.490 44.400 5.770 44.520 ;
        RECT 6.620 44.400 11.520 44.520 ;
        RECT 12.370 44.400 17.270 44.520 ;
        RECT 18.120 44.400 23.020 44.520 ;
        RECT 23.870 44.400 28.770 44.520 ;
        RECT 29.620 44.400 34.520 44.520 ;
        RECT 35.370 44.400 40.270 44.520 ;
        RECT 41.120 44.400 46.020 44.520 ;
        RECT 46.870 44.400 51.770 44.520 ;
        RECT 52.620 44.400 57.520 44.520 ;
        RECT 58.370 44.400 63.270 44.520 ;
        RECT 64.120 44.400 69.020 44.520 ;
        RECT 69.870 44.400 74.770 44.520 ;
        RECT 75.620 44.400 80.520 44.520 ;
        RECT 81.370 44.400 86.270 44.520 ;
        RECT 87.120 44.400 92.020 44.520 ;
        RECT 92.870 44.400 146.400 44.520 ;
        RECT -45.490 42.370 146.400 44.400 ;
        RECT -45.490 42.250 4.160 42.370 ;
        RECT 5.010 42.250 9.910 42.370 ;
        RECT 10.760 42.250 15.660 42.370 ;
        RECT 16.510 42.250 21.410 42.370 ;
        RECT 22.260 42.250 27.160 42.370 ;
        RECT 28.010 42.250 32.910 42.370 ;
        RECT 33.760 42.250 38.660 42.370 ;
        RECT 39.510 42.250 44.410 42.370 ;
        RECT 45.260 42.250 50.160 42.370 ;
        RECT 51.010 42.250 55.910 42.370 ;
        RECT 56.760 42.250 61.660 42.370 ;
        RECT 62.510 42.250 67.410 42.370 ;
        RECT 68.260 42.250 73.160 42.370 ;
        RECT 74.010 42.250 78.910 42.370 ;
        RECT 79.760 42.250 84.660 42.370 ;
        RECT 85.510 42.250 90.410 42.370 ;
        RECT 91.260 42.250 146.400 42.370 ;
        RECT 94.940 41.550 146.400 42.250 ;
        RECT -45.490 41.430 5.770 41.550 ;
        RECT 6.620 41.430 11.520 41.550 ;
        RECT 12.370 41.430 17.270 41.550 ;
        RECT 18.120 41.430 23.020 41.550 ;
        RECT 23.870 41.430 28.770 41.550 ;
        RECT 29.620 41.430 34.520 41.550 ;
        RECT 35.370 41.430 40.270 41.550 ;
        RECT 41.120 41.430 46.020 41.550 ;
        RECT 46.870 41.430 51.770 41.550 ;
        RECT 52.620 41.430 57.520 41.550 ;
        RECT 58.370 41.430 63.270 41.550 ;
        RECT 64.120 41.430 69.020 41.550 ;
        RECT 69.870 41.430 74.770 41.550 ;
        RECT 75.620 41.430 80.520 41.550 ;
        RECT 81.370 41.430 86.270 41.550 ;
        RECT 87.120 41.430 92.020 41.550 ;
        RECT 92.870 41.430 146.400 41.550 ;
        RECT -45.490 39.960 146.400 41.430 ;
        RECT -45.490 39.840 4.160 39.960 ;
        RECT 5.010 39.840 9.910 39.960 ;
        RECT 10.760 39.840 15.660 39.960 ;
        RECT 16.510 39.840 21.410 39.960 ;
        RECT 22.260 39.840 27.160 39.960 ;
        RECT 28.010 39.840 32.910 39.960 ;
        RECT 33.760 39.840 38.660 39.960 ;
        RECT 39.510 39.840 44.410 39.960 ;
        RECT 45.260 39.840 50.160 39.960 ;
        RECT 51.010 39.840 55.910 39.960 ;
        RECT 56.760 39.840 61.660 39.960 ;
        RECT 62.510 39.840 67.410 39.960 ;
        RECT 68.260 39.840 73.160 39.960 ;
        RECT 74.010 39.840 78.910 39.960 ;
        RECT 79.760 39.840 84.660 39.960 ;
        RECT 85.510 39.840 90.410 39.960 ;
        RECT 91.260 39.840 146.400 39.960 ;
        RECT 94.940 39.140 146.400 39.840 ;
        RECT -45.490 39.020 5.770 39.140 ;
        RECT 6.620 39.020 11.520 39.140 ;
        RECT 12.370 39.020 17.270 39.140 ;
        RECT 18.120 39.020 23.020 39.140 ;
        RECT 23.870 39.020 28.770 39.140 ;
        RECT 29.620 39.020 34.520 39.140 ;
        RECT 35.370 39.020 40.270 39.140 ;
        RECT 41.120 39.020 46.020 39.140 ;
        RECT 46.870 39.020 51.770 39.140 ;
        RECT 52.620 39.020 57.520 39.140 ;
        RECT 58.370 39.020 63.270 39.140 ;
        RECT 64.120 39.020 69.020 39.140 ;
        RECT 69.870 39.020 74.770 39.140 ;
        RECT 75.620 39.020 80.520 39.140 ;
        RECT 81.370 39.020 86.270 39.140 ;
        RECT 87.120 39.020 92.020 39.140 ;
        RECT 92.870 39.020 146.400 39.140 ;
        RECT -45.490 37.900 146.400 39.020 ;
        RECT -45.490 37.830 2.180 37.900 ;
        RECT 3.040 37.830 7.930 37.900 ;
        RECT 8.790 37.830 13.680 37.900 ;
        RECT 14.540 37.830 19.430 37.900 ;
        RECT 20.290 37.830 25.180 37.900 ;
        RECT 26.040 37.830 30.930 37.900 ;
        RECT 31.790 37.830 36.680 37.900 ;
        RECT 37.540 37.830 42.430 37.900 ;
        RECT 43.290 37.830 48.180 37.900 ;
        RECT 49.040 37.830 53.930 37.900 ;
        RECT 54.790 37.830 59.680 37.900 ;
        RECT 60.540 37.830 65.430 37.900 ;
        RECT 66.290 37.830 71.180 37.900 ;
        RECT 72.040 37.830 76.930 37.900 ;
        RECT 77.790 37.830 82.680 37.900 ;
        RECT 83.540 37.830 88.430 37.900 ;
        RECT 89.290 37.830 146.400 37.900 ;
        RECT 94.940 36.320 146.400 37.830 ;
        RECT -45.490 36.230 7.730 36.320 ;
        RECT 8.590 36.230 13.480 36.320 ;
        RECT 14.340 36.230 19.230 36.320 ;
        RECT 20.090 36.230 24.980 36.320 ;
        RECT 25.840 36.230 30.730 36.320 ;
        RECT 31.590 36.230 36.480 36.320 ;
        RECT 37.340 36.230 42.230 36.320 ;
        RECT 43.090 36.230 47.980 36.320 ;
        RECT 48.840 36.230 53.730 36.320 ;
        RECT 54.590 36.230 59.480 36.320 ;
        RECT 60.340 36.230 65.230 36.320 ;
        RECT 66.090 36.230 70.980 36.320 ;
        RECT 71.840 36.230 76.730 36.320 ;
        RECT 77.590 36.230 82.480 36.320 ;
        RECT 83.340 36.230 88.230 36.320 ;
        RECT 89.090 36.230 93.980 36.320 ;
        RECT 94.840 36.230 146.400 36.320 ;
        RECT -45.490 35.490 146.400 36.230 ;
        RECT -45.490 35.420 2.180 35.490 ;
        RECT 3.040 35.420 7.930 35.490 ;
        RECT 8.790 35.420 13.680 35.490 ;
        RECT 14.540 35.420 19.430 35.490 ;
        RECT 20.290 35.420 25.180 35.490 ;
        RECT 26.040 35.420 30.930 35.490 ;
        RECT 31.790 35.420 36.680 35.490 ;
        RECT 37.540 35.420 42.430 35.490 ;
        RECT 43.290 35.420 48.180 35.490 ;
        RECT 49.040 35.420 53.930 35.490 ;
        RECT 54.790 35.420 59.680 35.490 ;
        RECT 60.540 35.420 65.430 35.490 ;
        RECT 66.290 35.420 71.180 35.490 ;
        RECT 72.040 35.420 76.930 35.490 ;
        RECT 77.790 35.420 82.680 35.490 ;
        RECT 83.540 35.420 88.430 35.490 ;
        RECT 89.290 35.420 146.400 35.490 ;
        RECT 94.940 33.910 146.400 35.420 ;
        RECT -45.490 33.820 7.730 33.910 ;
        RECT 8.590 33.820 13.480 33.910 ;
        RECT 14.340 33.820 19.230 33.910 ;
        RECT 20.090 33.820 24.980 33.910 ;
        RECT 25.840 33.820 30.730 33.910 ;
        RECT 31.590 33.820 36.480 33.910 ;
        RECT 37.340 33.820 42.230 33.910 ;
        RECT 43.090 33.820 47.980 33.910 ;
        RECT 48.840 33.820 53.730 33.910 ;
        RECT 54.590 33.820 59.480 33.910 ;
        RECT 60.340 33.820 65.230 33.910 ;
        RECT 66.090 33.820 70.980 33.910 ;
        RECT 71.840 33.820 76.730 33.910 ;
        RECT 77.590 33.820 82.480 33.910 ;
        RECT 83.340 33.820 88.230 33.910 ;
        RECT 89.090 33.820 93.980 33.910 ;
        RECT 94.840 33.820 146.400 33.910 ;
        RECT -45.490 33.080 146.400 33.820 ;
        RECT -45.490 33.010 2.180 33.080 ;
        RECT 3.040 33.010 7.930 33.080 ;
        RECT 8.790 33.010 13.680 33.080 ;
        RECT 14.540 33.010 19.430 33.080 ;
        RECT 20.290 33.010 25.180 33.080 ;
        RECT 26.040 33.010 30.930 33.080 ;
        RECT 31.790 33.010 36.680 33.080 ;
        RECT 37.540 33.010 42.430 33.080 ;
        RECT 43.290 33.010 48.180 33.080 ;
        RECT 49.040 33.010 53.930 33.080 ;
        RECT 54.790 33.010 59.680 33.080 ;
        RECT 60.540 33.010 65.430 33.080 ;
        RECT 66.290 33.010 71.180 33.080 ;
        RECT 72.040 33.010 76.930 33.080 ;
        RECT 77.790 33.010 82.680 33.080 ;
        RECT 83.540 33.010 88.430 33.080 ;
        RECT 89.290 33.010 146.400 33.080 ;
        RECT 94.940 31.500 146.400 33.010 ;
        RECT -45.490 31.410 7.730 31.500 ;
        RECT 8.590 31.410 13.480 31.500 ;
        RECT 14.340 31.410 19.230 31.500 ;
        RECT 20.090 31.410 24.980 31.500 ;
        RECT 25.840 31.410 30.730 31.500 ;
        RECT 31.590 31.410 36.480 31.500 ;
        RECT 37.340 31.410 42.230 31.500 ;
        RECT 43.090 31.410 47.980 31.500 ;
        RECT 48.840 31.410 53.730 31.500 ;
        RECT 54.590 31.410 59.480 31.500 ;
        RECT 60.340 31.410 65.230 31.500 ;
        RECT 66.090 31.410 70.980 31.500 ;
        RECT 71.840 31.410 76.730 31.500 ;
        RECT 77.590 31.410 82.480 31.500 ;
        RECT 83.340 31.410 88.230 31.500 ;
        RECT 89.090 31.410 93.980 31.500 ;
        RECT 94.840 31.410 146.400 31.500 ;
        RECT -45.490 30.670 146.400 31.410 ;
        RECT -45.490 30.600 2.180 30.670 ;
        RECT 3.040 30.600 7.930 30.670 ;
        RECT 8.790 30.600 13.680 30.670 ;
        RECT 14.540 30.600 19.430 30.670 ;
        RECT 20.290 30.600 25.180 30.670 ;
        RECT 26.040 30.600 30.930 30.670 ;
        RECT 31.790 30.600 36.680 30.670 ;
        RECT 37.540 30.600 42.430 30.670 ;
        RECT 43.290 30.600 48.180 30.670 ;
        RECT 49.040 30.600 53.930 30.670 ;
        RECT 54.790 30.600 59.680 30.670 ;
        RECT 60.540 30.600 65.430 30.670 ;
        RECT 66.290 30.600 71.180 30.670 ;
        RECT 72.040 30.600 76.930 30.670 ;
        RECT 77.790 30.600 82.680 30.670 ;
        RECT 83.540 30.600 88.430 30.670 ;
        RECT 89.290 30.600 146.400 30.670 ;
        RECT 94.940 29.090 146.400 30.600 ;
        RECT -45.490 29.000 7.730 29.090 ;
        RECT 8.590 29.000 13.480 29.090 ;
        RECT 14.340 29.000 19.230 29.090 ;
        RECT 20.090 29.000 24.980 29.090 ;
        RECT 25.840 29.000 30.730 29.090 ;
        RECT 31.590 29.000 36.480 29.090 ;
        RECT 37.340 29.000 42.230 29.090 ;
        RECT 43.090 29.000 47.980 29.090 ;
        RECT 48.840 29.000 53.730 29.090 ;
        RECT 54.590 29.000 59.480 29.090 ;
        RECT 60.340 29.000 65.230 29.090 ;
        RECT 66.090 29.000 70.980 29.090 ;
        RECT 71.840 29.000 76.730 29.090 ;
        RECT 77.590 29.000 82.480 29.090 ;
        RECT 83.340 29.000 88.230 29.090 ;
        RECT 89.090 29.000 93.980 29.090 ;
        RECT 94.840 29.000 146.400 29.090 ;
        RECT -45.490 27.850 146.400 29.000 ;
        RECT -45.490 27.790 2.180 27.850 ;
        RECT 3.040 27.790 7.930 27.850 ;
        RECT 8.790 27.790 13.680 27.850 ;
        RECT 14.540 27.790 19.430 27.850 ;
        RECT 20.290 27.790 25.180 27.850 ;
        RECT 26.040 27.790 30.930 27.850 ;
        RECT 31.790 27.790 36.680 27.850 ;
        RECT 37.540 27.790 42.430 27.850 ;
        RECT 43.290 27.790 48.180 27.850 ;
        RECT 49.040 27.790 53.930 27.850 ;
        RECT 54.790 27.790 59.680 27.850 ;
        RECT 60.540 27.790 65.430 27.850 ;
        RECT 66.290 27.790 71.180 27.850 ;
        RECT 72.040 27.790 76.930 27.850 ;
        RECT 77.790 27.790 82.680 27.850 ;
        RECT 83.540 27.790 88.430 27.850 ;
        RECT 89.290 27.790 146.400 27.850 ;
        RECT 94.940 26.280 146.400 27.790 ;
        RECT -45.490 26.190 7.730 26.280 ;
        RECT 8.590 26.190 13.480 26.280 ;
        RECT 14.340 26.190 19.230 26.280 ;
        RECT 20.090 26.190 24.980 26.280 ;
        RECT 25.840 26.190 30.730 26.280 ;
        RECT 31.590 26.190 36.480 26.280 ;
        RECT 37.340 26.190 42.230 26.280 ;
        RECT 43.090 26.190 47.980 26.280 ;
        RECT 48.840 26.190 53.730 26.280 ;
        RECT 54.590 26.190 59.480 26.280 ;
        RECT 60.340 26.190 65.230 26.280 ;
        RECT 66.090 26.190 70.980 26.280 ;
        RECT 71.840 26.190 76.730 26.280 ;
        RECT 77.590 26.190 82.480 26.280 ;
        RECT 83.340 26.190 88.230 26.280 ;
        RECT 89.090 26.190 93.980 26.280 ;
        RECT 94.840 26.190 146.400 26.280 ;
        RECT -45.490 25.450 146.400 26.190 ;
        RECT -45.490 25.380 2.180 25.450 ;
        RECT 3.040 25.380 7.930 25.450 ;
        RECT 8.790 25.380 13.680 25.450 ;
        RECT 14.540 25.380 19.430 25.450 ;
        RECT 20.290 25.380 25.180 25.450 ;
        RECT 26.040 25.380 30.930 25.450 ;
        RECT 31.790 25.380 36.680 25.450 ;
        RECT 37.540 25.380 42.430 25.450 ;
        RECT 43.290 25.380 48.180 25.450 ;
        RECT 49.040 25.380 53.930 25.450 ;
        RECT 54.790 25.380 59.680 25.450 ;
        RECT 60.540 25.380 65.430 25.450 ;
        RECT 66.290 25.380 71.180 25.450 ;
        RECT 72.040 25.380 76.930 25.450 ;
        RECT 77.790 25.380 82.680 25.450 ;
        RECT 83.540 25.380 88.430 25.450 ;
        RECT 89.290 25.380 146.400 25.450 ;
        RECT 94.940 23.870 146.400 25.380 ;
        RECT -45.490 23.780 7.730 23.870 ;
        RECT 8.590 23.780 13.480 23.870 ;
        RECT 14.340 23.780 19.230 23.870 ;
        RECT 20.090 23.780 24.980 23.870 ;
        RECT 25.840 23.780 30.730 23.870 ;
        RECT 31.590 23.780 36.480 23.870 ;
        RECT 37.340 23.780 42.230 23.870 ;
        RECT 43.090 23.780 47.980 23.870 ;
        RECT 48.840 23.780 53.730 23.870 ;
        RECT 54.590 23.780 59.480 23.870 ;
        RECT 60.340 23.780 65.230 23.870 ;
        RECT 66.090 23.780 70.980 23.870 ;
        RECT 71.840 23.780 76.730 23.870 ;
        RECT 77.590 23.780 82.480 23.870 ;
        RECT 83.340 23.780 88.230 23.870 ;
        RECT 89.090 23.780 93.980 23.870 ;
        RECT 94.840 23.780 146.400 23.870 ;
        RECT -45.490 23.040 146.400 23.780 ;
        RECT -45.490 22.970 2.180 23.040 ;
        RECT 3.040 22.970 7.930 23.040 ;
        RECT 8.790 22.970 13.680 23.040 ;
        RECT 14.540 22.970 19.430 23.040 ;
        RECT 20.290 22.970 25.180 23.040 ;
        RECT 26.040 22.970 30.930 23.040 ;
        RECT 31.790 22.970 36.680 23.040 ;
        RECT 37.540 22.970 42.430 23.040 ;
        RECT 43.290 22.970 48.180 23.040 ;
        RECT 49.040 22.970 53.930 23.040 ;
        RECT 54.790 22.970 59.680 23.040 ;
        RECT 60.540 22.970 65.430 23.040 ;
        RECT 66.290 22.970 71.180 23.040 ;
        RECT 72.040 22.970 76.930 23.040 ;
        RECT 77.790 22.970 82.680 23.040 ;
        RECT 83.540 22.970 88.430 23.040 ;
        RECT 89.290 22.970 146.400 23.040 ;
        RECT 94.940 21.460 146.400 22.970 ;
        RECT -45.490 21.370 7.730 21.460 ;
        RECT 8.590 21.370 13.480 21.460 ;
        RECT 14.340 21.370 19.230 21.460 ;
        RECT 20.090 21.370 24.980 21.460 ;
        RECT 25.840 21.370 30.730 21.460 ;
        RECT 31.590 21.370 36.480 21.460 ;
        RECT 37.340 21.370 42.230 21.460 ;
        RECT 43.090 21.370 47.980 21.460 ;
        RECT 48.840 21.370 53.730 21.460 ;
        RECT 54.590 21.370 59.480 21.460 ;
        RECT 60.340 21.370 65.230 21.460 ;
        RECT 66.090 21.370 70.980 21.460 ;
        RECT 71.840 21.370 76.730 21.460 ;
        RECT 77.590 21.370 82.480 21.460 ;
        RECT 83.340 21.370 88.230 21.460 ;
        RECT 89.090 21.370 93.980 21.460 ;
        RECT 94.840 21.370 146.400 21.460 ;
        RECT -45.490 20.630 146.400 21.370 ;
        RECT -45.490 20.560 2.180 20.630 ;
        RECT 3.040 20.560 7.930 20.630 ;
        RECT 8.790 20.560 13.680 20.630 ;
        RECT 14.540 20.560 19.430 20.630 ;
        RECT 20.290 20.560 25.180 20.630 ;
        RECT 26.040 20.560 30.930 20.630 ;
        RECT 31.790 20.560 36.680 20.630 ;
        RECT 37.540 20.560 42.430 20.630 ;
        RECT 43.290 20.560 48.180 20.630 ;
        RECT 49.040 20.560 53.930 20.630 ;
        RECT 54.790 20.560 59.680 20.630 ;
        RECT 60.540 20.560 65.430 20.630 ;
        RECT 66.290 20.560 71.180 20.630 ;
        RECT 72.040 20.560 76.930 20.630 ;
        RECT 77.790 20.560 82.680 20.630 ;
        RECT 83.540 20.560 88.430 20.630 ;
        RECT 89.290 20.560 146.400 20.630 ;
        RECT 94.940 19.050 146.400 20.560 ;
        RECT -45.490 18.960 7.730 19.050 ;
        RECT 8.590 18.960 13.480 19.050 ;
        RECT 14.340 18.960 19.230 19.050 ;
        RECT 20.090 18.960 24.980 19.050 ;
        RECT 25.840 18.960 30.730 19.050 ;
        RECT 31.590 18.960 36.480 19.050 ;
        RECT 37.340 18.960 42.230 19.050 ;
        RECT 43.090 18.960 47.980 19.050 ;
        RECT 48.840 18.960 53.730 19.050 ;
        RECT 54.590 18.960 59.480 19.050 ;
        RECT 60.340 18.960 65.230 19.050 ;
        RECT 66.090 18.960 70.980 19.050 ;
        RECT 71.840 18.960 76.730 19.050 ;
        RECT 77.590 18.960 82.480 19.050 ;
        RECT 83.340 18.960 88.230 19.050 ;
        RECT 89.090 18.960 93.980 19.050 ;
        RECT 94.840 18.960 146.400 19.050 ;
        RECT -45.490 18.220 146.400 18.960 ;
        RECT -45.490 18.150 2.180 18.220 ;
        RECT 3.040 18.150 7.930 18.220 ;
        RECT 8.790 18.150 13.680 18.220 ;
        RECT 14.540 18.150 19.430 18.220 ;
        RECT 20.290 18.150 25.180 18.220 ;
        RECT 26.040 18.150 30.930 18.220 ;
        RECT 31.790 18.150 36.680 18.220 ;
        RECT 37.540 18.150 42.430 18.220 ;
        RECT 43.290 18.150 48.180 18.220 ;
        RECT 49.040 18.150 53.930 18.220 ;
        RECT 54.790 18.150 59.680 18.220 ;
        RECT 60.540 18.150 65.430 18.220 ;
        RECT 66.290 18.150 71.180 18.220 ;
        RECT 72.040 18.150 76.930 18.220 ;
        RECT 77.790 18.150 82.680 18.220 ;
        RECT 83.540 18.150 88.430 18.220 ;
        RECT 89.290 18.150 146.400 18.220 ;
        RECT 94.940 16.640 146.400 18.150 ;
        RECT -45.490 16.550 7.730 16.640 ;
        RECT 8.590 16.550 13.480 16.640 ;
        RECT 14.340 16.550 19.230 16.640 ;
        RECT 20.090 16.550 24.980 16.640 ;
        RECT 25.840 16.550 30.730 16.640 ;
        RECT 31.590 16.550 36.480 16.640 ;
        RECT 37.340 16.550 42.230 16.640 ;
        RECT 43.090 16.550 47.980 16.640 ;
        RECT 48.840 16.550 53.730 16.640 ;
        RECT 54.590 16.550 59.480 16.640 ;
        RECT 60.340 16.550 65.230 16.640 ;
        RECT 66.090 16.550 70.980 16.640 ;
        RECT 71.840 16.550 76.730 16.640 ;
        RECT 77.590 16.550 82.480 16.640 ;
        RECT 83.340 16.550 88.230 16.640 ;
        RECT 89.090 16.550 93.980 16.640 ;
        RECT 94.840 16.550 146.400 16.640 ;
        RECT -45.490 15.810 146.400 16.550 ;
        RECT -45.490 15.740 2.180 15.810 ;
        RECT 3.040 15.740 7.930 15.810 ;
        RECT 8.790 15.740 13.680 15.810 ;
        RECT 14.540 15.740 19.430 15.810 ;
        RECT 20.290 15.740 25.180 15.810 ;
        RECT 26.040 15.740 30.930 15.810 ;
        RECT 31.790 15.740 36.680 15.810 ;
        RECT 37.540 15.740 42.430 15.810 ;
        RECT 43.290 15.740 48.180 15.810 ;
        RECT 49.040 15.740 53.930 15.810 ;
        RECT 54.790 15.740 59.680 15.810 ;
        RECT 60.540 15.740 65.430 15.810 ;
        RECT 66.290 15.740 71.180 15.810 ;
        RECT 72.040 15.740 76.930 15.810 ;
        RECT 77.790 15.740 82.680 15.810 ;
        RECT 83.540 15.740 88.430 15.810 ;
        RECT 89.290 15.740 146.400 15.810 ;
        RECT 94.940 14.230 146.400 15.740 ;
        RECT -45.490 14.140 7.730 14.230 ;
        RECT 8.590 14.140 13.480 14.230 ;
        RECT 14.340 14.140 19.230 14.230 ;
        RECT 20.090 14.140 24.980 14.230 ;
        RECT 25.840 14.140 30.730 14.230 ;
        RECT 31.590 14.140 36.480 14.230 ;
        RECT 37.340 14.140 42.230 14.230 ;
        RECT 43.090 14.140 47.980 14.230 ;
        RECT 48.840 14.140 53.730 14.230 ;
        RECT 54.590 14.140 59.480 14.230 ;
        RECT 60.340 14.140 65.230 14.230 ;
        RECT 66.090 14.140 70.980 14.230 ;
        RECT 71.840 14.140 76.730 14.230 ;
        RECT 77.590 14.140 82.480 14.230 ;
        RECT 83.340 14.140 88.230 14.230 ;
        RECT 89.090 14.140 93.980 14.230 ;
        RECT 94.840 14.140 146.400 14.230 ;
        RECT -45.490 13.400 146.400 14.140 ;
        RECT -45.490 13.330 2.180 13.400 ;
        RECT 3.040 13.330 7.930 13.400 ;
        RECT 8.790 13.330 13.680 13.400 ;
        RECT 14.540 13.330 19.430 13.400 ;
        RECT 20.290 13.330 25.180 13.400 ;
        RECT 26.040 13.330 30.930 13.400 ;
        RECT 31.790 13.330 36.680 13.400 ;
        RECT 37.540 13.330 42.430 13.400 ;
        RECT 43.290 13.330 48.180 13.400 ;
        RECT 49.040 13.330 53.930 13.400 ;
        RECT 54.790 13.330 59.680 13.400 ;
        RECT 60.540 13.330 65.430 13.400 ;
        RECT 66.290 13.330 71.180 13.400 ;
        RECT 72.040 13.330 76.930 13.400 ;
        RECT 77.790 13.330 82.680 13.400 ;
        RECT 83.540 13.330 88.430 13.400 ;
        RECT 89.290 13.330 146.400 13.400 ;
        RECT 94.940 11.820 146.400 13.330 ;
        RECT -45.490 11.730 7.730 11.820 ;
        RECT 8.590 11.730 13.480 11.820 ;
        RECT 14.340 11.730 19.230 11.820 ;
        RECT 20.090 11.730 24.980 11.820 ;
        RECT 25.840 11.730 30.730 11.820 ;
        RECT 31.590 11.730 36.480 11.820 ;
        RECT 37.340 11.730 42.230 11.820 ;
        RECT 43.090 11.730 47.980 11.820 ;
        RECT 48.840 11.730 53.730 11.820 ;
        RECT 54.590 11.730 59.480 11.820 ;
        RECT 60.340 11.730 65.230 11.820 ;
        RECT 66.090 11.730 70.980 11.820 ;
        RECT 71.840 11.730 76.730 11.820 ;
        RECT 77.590 11.730 82.480 11.820 ;
        RECT 83.340 11.730 88.230 11.820 ;
        RECT 89.090 11.730 93.980 11.820 ;
        RECT 94.840 11.730 146.400 11.820 ;
        RECT -45.490 10.990 146.400 11.730 ;
        RECT -45.490 10.920 2.180 10.990 ;
        RECT 3.040 10.920 7.930 10.990 ;
        RECT 8.790 10.920 13.680 10.990 ;
        RECT 14.540 10.920 19.430 10.990 ;
        RECT 20.290 10.920 25.180 10.990 ;
        RECT 26.040 10.920 30.930 10.990 ;
        RECT 31.790 10.920 36.680 10.990 ;
        RECT 37.540 10.920 42.430 10.990 ;
        RECT 43.290 10.920 48.180 10.990 ;
        RECT 49.040 10.920 53.930 10.990 ;
        RECT 54.790 10.920 59.680 10.990 ;
        RECT 60.540 10.920 65.430 10.990 ;
        RECT 66.290 10.920 71.180 10.990 ;
        RECT 72.040 10.920 76.930 10.990 ;
        RECT 77.790 10.920 82.680 10.990 ;
        RECT 83.540 10.920 88.430 10.990 ;
        RECT 89.290 10.920 146.400 10.990 ;
        RECT 94.940 9.410 146.400 10.920 ;
        RECT -45.490 9.320 7.730 9.410 ;
        RECT 8.590 9.320 13.480 9.410 ;
        RECT 14.340 9.320 19.230 9.410 ;
        RECT 20.090 9.320 24.980 9.410 ;
        RECT 25.840 9.320 30.730 9.410 ;
        RECT 31.590 9.320 36.480 9.410 ;
        RECT 37.340 9.320 42.230 9.410 ;
        RECT 43.090 9.320 47.980 9.410 ;
        RECT 48.840 9.320 53.730 9.410 ;
        RECT 54.590 9.320 59.480 9.410 ;
        RECT 60.340 9.320 65.230 9.410 ;
        RECT 66.090 9.320 70.980 9.410 ;
        RECT 71.840 9.320 76.730 9.410 ;
        RECT 77.590 9.320 82.480 9.410 ;
        RECT 83.340 9.320 88.230 9.410 ;
        RECT 89.090 9.320 93.980 9.410 ;
        RECT 94.840 9.320 146.400 9.410 ;
        RECT -45.490 8.160 146.400 9.320 ;
        RECT -45.490 8.100 2.180 8.160 ;
        RECT 3.040 8.100 7.930 8.160 ;
        RECT 8.790 8.100 13.680 8.160 ;
        RECT 14.540 8.100 19.430 8.160 ;
        RECT 20.290 8.100 25.180 8.160 ;
        RECT 26.040 8.100 30.930 8.160 ;
        RECT 31.790 8.100 36.680 8.160 ;
        RECT 37.540 8.100 42.430 8.160 ;
        RECT 43.290 8.100 48.180 8.160 ;
        RECT 49.040 8.100 53.930 8.160 ;
        RECT 54.790 8.100 59.680 8.160 ;
        RECT 60.540 8.100 65.430 8.160 ;
        RECT 66.290 8.100 71.180 8.160 ;
        RECT 72.040 8.100 76.930 8.160 ;
        RECT 77.790 8.100 82.680 8.160 ;
        RECT 83.540 8.100 88.430 8.160 ;
        RECT 89.290 8.100 146.400 8.160 ;
        RECT 94.940 6.590 146.400 8.100 ;
        RECT -45.490 6.500 7.730 6.590 ;
        RECT 8.590 6.500 13.480 6.590 ;
        RECT 14.340 6.500 19.230 6.590 ;
        RECT 20.090 6.500 24.980 6.590 ;
        RECT 25.840 6.500 30.730 6.590 ;
        RECT 31.590 6.500 36.480 6.590 ;
        RECT 37.340 6.500 42.230 6.590 ;
        RECT 43.090 6.500 47.980 6.590 ;
        RECT 48.840 6.500 53.730 6.590 ;
        RECT 54.590 6.500 59.480 6.590 ;
        RECT 60.340 6.500 65.230 6.590 ;
        RECT 66.090 6.500 70.980 6.590 ;
        RECT 71.840 6.500 76.730 6.590 ;
        RECT 77.590 6.500 82.480 6.590 ;
        RECT 83.340 6.500 88.230 6.590 ;
        RECT 89.090 6.500 93.980 6.590 ;
        RECT 94.840 6.500 146.400 6.590 ;
        RECT -45.490 5.760 146.400 6.500 ;
        RECT -45.490 5.690 2.180 5.760 ;
        RECT 3.040 5.690 7.930 5.760 ;
        RECT 8.790 5.690 13.680 5.760 ;
        RECT 14.540 5.690 19.430 5.760 ;
        RECT 20.290 5.690 25.180 5.760 ;
        RECT 26.040 5.690 30.930 5.760 ;
        RECT 31.790 5.690 36.680 5.760 ;
        RECT 37.540 5.690 42.430 5.760 ;
        RECT 43.290 5.690 48.180 5.760 ;
        RECT 49.040 5.690 53.930 5.760 ;
        RECT 54.790 5.690 59.680 5.760 ;
        RECT 60.540 5.690 65.430 5.760 ;
        RECT 66.290 5.690 71.180 5.760 ;
        RECT 72.040 5.690 76.930 5.760 ;
        RECT 77.790 5.690 82.680 5.760 ;
        RECT 83.540 5.690 88.430 5.760 ;
        RECT 89.290 5.690 146.400 5.760 ;
        RECT 94.940 4.180 146.400 5.690 ;
        RECT -45.490 4.090 7.730 4.180 ;
        RECT 8.590 4.090 13.480 4.180 ;
        RECT 14.340 4.090 19.230 4.180 ;
        RECT 20.090 4.090 24.980 4.180 ;
        RECT 25.840 4.090 30.730 4.180 ;
        RECT 31.590 4.090 36.480 4.180 ;
        RECT 37.340 4.090 42.230 4.180 ;
        RECT 43.090 4.090 47.980 4.180 ;
        RECT 48.840 4.090 53.730 4.180 ;
        RECT 54.590 4.090 59.480 4.180 ;
        RECT 60.340 4.090 65.230 4.180 ;
        RECT 66.090 4.090 70.980 4.180 ;
        RECT 71.840 4.090 76.730 4.180 ;
        RECT 77.590 4.090 82.480 4.180 ;
        RECT 83.340 4.090 88.230 4.180 ;
        RECT 89.090 4.090 93.980 4.180 ;
        RECT 94.840 4.090 146.400 4.180 ;
        RECT -45.490 3.350 146.400 4.090 ;
        RECT -45.490 3.280 2.180 3.350 ;
        RECT 3.040 3.280 7.930 3.350 ;
        RECT 8.790 3.280 13.680 3.350 ;
        RECT 14.540 3.280 19.430 3.350 ;
        RECT 20.290 3.280 25.180 3.350 ;
        RECT 26.040 3.280 30.930 3.350 ;
        RECT 31.790 3.280 36.680 3.350 ;
        RECT 37.540 3.280 42.430 3.350 ;
        RECT 43.290 3.280 48.180 3.350 ;
        RECT 49.040 3.280 53.930 3.350 ;
        RECT 54.790 3.280 59.680 3.350 ;
        RECT 60.540 3.280 65.430 3.350 ;
        RECT 66.290 3.280 71.180 3.350 ;
        RECT 72.040 3.280 76.930 3.350 ;
        RECT 77.790 3.280 82.680 3.350 ;
        RECT 83.540 3.280 88.430 3.350 ;
        RECT 89.290 3.280 146.400 3.350 ;
        RECT 94.940 1.770 146.400 3.280 ;
        RECT -45.490 1.680 7.730 1.770 ;
        RECT 8.590 1.680 13.480 1.770 ;
        RECT 14.340 1.680 19.230 1.770 ;
        RECT 20.090 1.680 24.980 1.770 ;
        RECT 25.840 1.680 30.730 1.770 ;
        RECT 31.590 1.680 36.480 1.770 ;
        RECT 37.340 1.680 42.230 1.770 ;
        RECT 43.090 1.680 47.980 1.770 ;
        RECT 48.840 1.680 53.730 1.770 ;
        RECT 54.590 1.680 59.480 1.770 ;
        RECT 60.340 1.680 65.230 1.770 ;
        RECT 66.090 1.680 70.980 1.770 ;
        RECT 71.840 1.680 76.730 1.770 ;
        RECT 77.590 1.680 82.480 1.770 ;
        RECT 83.340 1.680 88.230 1.770 ;
        RECT 89.090 1.680 93.980 1.770 ;
        RECT 94.840 1.680 146.400 1.770 ;
        RECT -45.490 0.940 146.400 1.680 ;
        RECT -45.490 0.870 2.180 0.940 ;
        RECT 3.040 0.870 7.930 0.940 ;
        RECT 8.790 0.870 13.680 0.940 ;
        RECT 14.540 0.870 19.430 0.940 ;
        RECT 20.290 0.870 25.180 0.940 ;
        RECT 26.040 0.870 30.930 0.940 ;
        RECT 31.790 0.870 36.680 0.940 ;
        RECT 37.540 0.870 42.430 0.940 ;
        RECT 43.290 0.870 48.180 0.940 ;
        RECT 49.040 0.870 53.930 0.940 ;
        RECT 54.790 0.870 59.680 0.940 ;
        RECT 60.540 0.870 65.430 0.940 ;
        RECT 66.290 0.870 71.180 0.940 ;
        RECT 72.040 0.870 76.930 0.940 ;
        RECT 77.790 0.870 82.680 0.940 ;
        RECT 83.540 0.870 88.430 0.940 ;
        RECT 89.290 0.870 146.400 0.940 ;
        RECT 94.940 -0.640 146.400 0.870 ;
        RECT -45.490 -0.730 7.730 -0.640 ;
        RECT 8.590 -0.730 13.480 -0.640 ;
        RECT 14.340 -0.730 19.230 -0.640 ;
        RECT 20.090 -0.730 24.980 -0.640 ;
        RECT 25.840 -0.730 30.730 -0.640 ;
        RECT 31.590 -0.730 36.480 -0.640 ;
        RECT 37.340 -0.730 42.230 -0.640 ;
        RECT 43.090 -0.730 47.980 -0.640 ;
        RECT 48.840 -0.730 53.730 -0.640 ;
        RECT 54.590 -0.730 59.480 -0.640 ;
        RECT 60.340 -0.730 65.230 -0.640 ;
        RECT 66.090 -0.730 70.980 -0.640 ;
        RECT 71.840 -0.730 76.730 -0.640 ;
        RECT 77.590 -0.730 82.480 -0.640 ;
        RECT 83.340 -0.730 88.230 -0.640 ;
        RECT 89.090 -0.730 93.980 -0.640 ;
        RECT 94.840 -0.730 146.400 -0.640 ;
        RECT -45.490 -1.820 146.400 -0.730 ;
        RECT -45.490 -1.940 4.160 -1.820 ;
        RECT 5.010 -1.940 9.910 -1.820 ;
        RECT 10.760 -1.940 15.660 -1.820 ;
        RECT 16.510 -1.940 21.410 -1.820 ;
        RECT 22.260 -1.940 27.160 -1.820 ;
        RECT 28.010 -1.940 32.910 -1.820 ;
        RECT 33.760 -1.940 38.660 -1.820 ;
        RECT 39.510 -1.940 44.410 -1.820 ;
        RECT 45.260 -1.940 50.160 -1.820 ;
        RECT 51.010 -1.940 55.910 -1.820 ;
        RECT 56.760 -1.940 61.660 -1.820 ;
        RECT 62.510 -1.940 67.410 -1.820 ;
        RECT 68.260 -1.940 73.160 -1.820 ;
        RECT 74.010 -1.940 78.910 -1.820 ;
        RECT 79.760 -1.940 84.660 -1.820 ;
        RECT 85.510 -1.940 90.410 -1.820 ;
        RECT 91.260 -1.940 146.400 -1.820 ;
        RECT 94.940 -2.640 146.400 -1.940 ;
        RECT -45.490 -2.760 5.770 -2.640 ;
        RECT 6.620 -2.760 11.520 -2.640 ;
        RECT 12.370 -2.760 17.270 -2.640 ;
        RECT 18.120 -2.760 23.020 -2.640 ;
        RECT 23.870 -2.760 28.770 -2.640 ;
        RECT 29.620 -2.760 34.520 -2.640 ;
        RECT 35.370 -2.760 40.270 -2.640 ;
        RECT 41.120 -2.760 46.020 -2.640 ;
        RECT 46.870 -2.760 51.770 -2.640 ;
        RECT 52.620 -2.760 57.520 -2.640 ;
        RECT 58.370 -2.760 63.270 -2.640 ;
        RECT 64.120 -2.760 69.020 -2.640 ;
        RECT 69.870 -2.760 74.770 -2.640 ;
        RECT 75.620 -2.760 80.520 -2.640 ;
        RECT 81.370 -2.760 86.270 -2.640 ;
        RECT 87.120 -2.760 92.020 -2.640 ;
        RECT 92.870 -2.760 146.400 -2.640 ;
        RECT -45.490 -4.230 146.400 -2.760 ;
        RECT -45.490 -4.350 4.160 -4.230 ;
        RECT 5.010 -4.350 9.910 -4.230 ;
        RECT 10.760 -4.350 15.660 -4.230 ;
        RECT 16.510 -4.350 21.410 -4.230 ;
        RECT 22.260 -4.350 27.160 -4.230 ;
        RECT 28.010 -4.350 32.910 -4.230 ;
        RECT 33.760 -4.350 38.660 -4.230 ;
        RECT 39.510 -4.350 44.410 -4.230 ;
        RECT 45.260 -4.350 50.160 -4.230 ;
        RECT 51.010 -4.350 55.910 -4.230 ;
        RECT 56.760 -4.350 61.660 -4.230 ;
        RECT 62.510 -4.350 67.410 -4.230 ;
        RECT 68.260 -4.350 73.160 -4.230 ;
        RECT 74.010 -4.350 78.910 -4.230 ;
        RECT 79.760 -4.350 84.660 -4.230 ;
        RECT 85.510 -4.350 90.410 -4.230 ;
        RECT 91.260 -4.350 146.400 -4.230 ;
        RECT 94.940 -5.050 146.400 -4.350 ;
        RECT -45.490 -5.170 5.770 -5.050 ;
        RECT 6.620 -5.170 11.520 -5.050 ;
        RECT 12.370 -5.170 17.270 -5.050 ;
        RECT 18.120 -5.170 23.020 -5.050 ;
        RECT 23.870 -5.170 28.770 -5.050 ;
        RECT 29.620 -5.170 34.520 -5.050 ;
        RECT 35.370 -5.170 40.270 -5.050 ;
        RECT 41.120 -5.170 46.020 -5.050 ;
        RECT 46.870 -5.170 51.770 -5.050 ;
        RECT 52.620 -5.170 57.520 -5.050 ;
        RECT 58.370 -5.170 63.270 -5.050 ;
        RECT 64.120 -5.170 69.020 -5.050 ;
        RECT 69.870 -5.170 74.770 -5.050 ;
        RECT 75.620 -5.170 80.520 -5.050 ;
        RECT 81.370 -5.170 86.270 -5.050 ;
        RECT 87.120 -5.170 92.020 -5.050 ;
        RECT 92.870 -5.170 146.400 -5.050 ;
        RECT -45.490 -7.230 146.400 -5.170 ;
        RECT -45.490 -7.350 4.160 -7.230 ;
        RECT 5.010 -7.350 9.910 -7.230 ;
        RECT 10.760 -7.350 15.660 -7.230 ;
        RECT 16.510 -7.350 21.410 -7.230 ;
        RECT 22.260 -7.350 27.160 -7.230 ;
        RECT 28.010 -7.350 32.910 -7.230 ;
        RECT 33.760 -7.350 38.660 -7.230 ;
        RECT 39.510 -7.350 44.410 -7.230 ;
        RECT 45.260 -7.350 50.160 -7.230 ;
        RECT 51.010 -7.350 55.910 -7.230 ;
        RECT 56.760 -7.350 61.660 -7.230 ;
        RECT 62.510 -7.350 67.410 -7.230 ;
        RECT 68.260 -7.350 73.160 -7.230 ;
        RECT 74.010 -7.350 78.910 -7.230 ;
        RECT 79.760 -7.350 84.660 -7.230 ;
        RECT 85.510 -7.350 90.410 -7.230 ;
        RECT 91.260 -7.350 146.400 -7.230 ;
        RECT 94.940 -8.050 146.400 -7.350 ;
        RECT -45.490 -8.170 5.770 -8.050 ;
        RECT 6.620 -8.170 11.520 -8.050 ;
        RECT 12.370 -8.170 17.270 -8.050 ;
        RECT 18.120 -8.170 23.020 -8.050 ;
        RECT 23.870 -8.170 28.770 -8.050 ;
        RECT 29.620 -8.170 34.520 -8.050 ;
        RECT 35.370 -8.170 40.270 -8.050 ;
        RECT 41.120 -8.170 46.020 -8.050 ;
        RECT 46.870 -8.170 51.770 -8.050 ;
        RECT 52.620 -8.170 57.520 -8.050 ;
        RECT 58.370 -8.170 63.270 -8.050 ;
        RECT 64.120 -8.170 69.020 -8.050 ;
        RECT 69.870 -8.170 74.770 -8.050 ;
        RECT 75.620 -8.170 80.520 -8.050 ;
        RECT 81.370 -8.170 86.270 -8.050 ;
        RECT 87.120 -8.170 92.020 -8.050 ;
        RECT 92.870 -8.170 146.400 -8.050 ;
        RECT -45.490 -9.640 146.400 -8.170 ;
        RECT -45.490 -9.760 4.160 -9.640 ;
        RECT 5.010 -9.760 9.910 -9.640 ;
        RECT 10.760 -9.760 15.660 -9.640 ;
        RECT 16.510 -9.760 21.410 -9.640 ;
        RECT 22.260 -9.760 27.160 -9.640 ;
        RECT 28.010 -9.760 32.910 -9.640 ;
        RECT 33.760 -9.760 38.660 -9.640 ;
        RECT 39.510 -9.760 44.410 -9.640 ;
        RECT 45.260 -9.760 50.160 -9.640 ;
        RECT 51.010 -9.760 55.910 -9.640 ;
        RECT 56.760 -9.760 61.660 -9.640 ;
        RECT 62.510 -9.760 67.410 -9.640 ;
        RECT 68.260 -9.760 73.160 -9.640 ;
        RECT 74.010 -9.760 78.910 -9.640 ;
        RECT 79.760 -9.760 84.660 -9.640 ;
        RECT 85.510 -9.760 90.410 -9.640 ;
        RECT 91.260 -9.760 146.400 -9.640 ;
        RECT 94.940 -10.460 146.400 -9.760 ;
        RECT -45.490 -10.580 5.770 -10.460 ;
        RECT 6.620 -10.580 11.520 -10.460 ;
        RECT 12.370 -10.580 17.270 -10.460 ;
        RECT 18.120 -10.580 23.020 -10.460 ;
        RECT 23.870 -10.580 28.770 -10.460 ;
        RECT 29.620 -10.580 34.520 -10.460 ;
        RECT 35.370 -10.580 40.270 -10.460 ;
        RECT 41.120 -10.580 46.020 -10.460 ;
        RECT 46.870 -10.580 51.770 -10.460 ;
        RECT 52.620 -10.580 57.520 -10.460 ;
        RECT 58.370 -10.580 63.270 -10.460 ;
        RECT 64.120 -10.580 69.020 -10.460 ;
        RECT 69.870 -10.580 74.770 -10.460 ;
        RECT 75.620 -10.580 80.520 -10.460 ;
        RECT 81.370 -10.580 86.270 -10.460 ;
        RECT 87.120 -10.580 92.020 -10.460 ;
        RECT 92.870 -10.580 146.400 -10.460 ;
        RECT -45.490 -19.160 146.400 -10.580 ;
        RECT -45.490 -19.220 3.990 -19.160 ;
        RECT 4.880 -19.220 5.870 -19.160 ;
        RECT 6.760 -19.220 9.740 -19.160 ;
        RECT 10.630 -19.220 11.620 -19.160 ;
        RECT 12.510 -19.220 15.490 -19.160 ;
        RECT 16.380 -19.220 17.370 -19.160 ;
        RECT 18.260 -19.220 21.240 -19.160 ;
        RECT 22.130 -19.220 23.120 -19.160 ;
        RECT 24.010 -19.220 26.990 -19.160 ;
        RECT 27.880 -19.220 28.870 -19.160 ;
        RECT 29.760 -19.220 32.740 -19.160 ;
        RECT 33.630 -19.220 34.620 -19.160 ;
        RECT 35.510 -19.220 38.490 -19.160 ;
        RECT 39.380 -19.220 40.370 -19.160 ;
        RECT 41.260 -19.220 44.240 -19.160 ;
        RECT 45.130 -19.220 46.120 -19.160 ;
        RECT 47.010 -19.220 49.990 -19.160 ;
        RECT 50.880 -19.220 51.870 -19.160 ;
        RECT 52.760 -19.220 55.740 -19.160 ;
        RECT 56.630 -19.220 57.620 -19.160 ;
        RECT 58.510 -19.220 61.490 -19.160 ;
        RECT 62.380 -19.220 63.370 -19.160 ;
        RECT 64.260 -19.220 67.240 -19.160 ;
        RECT 68.130 -19.220 69.120 -19.160 ;
        RECT 70.010 -19.220 72.990 -19.160 ;
        RECT 73.880 -19.220 74.870 -19.160 ;
        RECT 75.760 -19.220 78.740 -19.160 ;
        RECT 79.630 -19.220 80.620 -19.160 ;
        RECT 81.510 -19.220 84.490 -19.160 ;
        RECT 85.380 -19.220 86.370 -19.160 ;
        RECT 87.260 -19.220 90.240 -19.160 ;
        RECT 91.130 -19.220 92.120 -19.160 ;
        RECT 93.010 -19.220 146.400 -19.160 ;
        RECT 94.940 -19.920 146.400 -19.220 ;
        RECT -45.490 -19.970 3.990 -19.920 ;
        RECT 4.880 -19.970 5.870 -19.920 ;
        RECT 6.760 -19.970 9.740 -19.920 ;
        RECT 10.630 -19.970 11.620 -19.920 ;
        RECT 12.510 -19.970 15.490 -19.920 ;
        RECT 16.380 -19.970 17.370 -19.920 ;
        RECT 18.260 -19.970 21.240 -19.920 ;
        RECT 22.130 -19.970 23.120 -19.920 ;
        RECT 24.010 -19.970 26.990 -19.920 ;
        RECT 27.880 -19.970 28.870 -19.920 ;
        RECT 29.760 -19.970 32.740 -19.920 ;
        RECT 33.630 -19.970 34.620 -19.920 ;
        RECT 35.510 -19.970 38.490 -19.920 ;
        RECT 39.380 -19.970 40.370 -19.920 ;
        RECT 41.260 -19.970 44.240 -19.920 ;
        RECT 45.130 -19.970 46.120 -19.920 ;
        RECT 47.010 -19.970 49.990 -19.920 ;
        RECT 50.880 -19.970 51.870 -19.920 ;
        RECT 52.760 -19.970 55.740 -19.920 ;
        RECT 56.630 -19.970 57.620 -19.920 ;
        RECT 58.510 -19.970 61.490 -19.920 ;
        RECT 62.380 -19.970 63.370 -19.920 ;
        RECT 64.260 -19.970 67.240 -19.920 ;
        RECT 68.130 -19.970 69.120 -19.920 ;
        RECT 70.010 -19.970 72.990 -19.920 ;
        RECT 73.880 -19.970 74.870 -19.920 ;
        RECT 75.760 -19.970 78.740 -19.920 ;
        RECT 79.630 -19.970 80.620 -19.920 ;
        RECT 81.510 -19.970 84.490 -19.920 ;
        RECT 85.380 -19.970 86.370 -19.920 ;
        RECT 87.260 -19.970 90.240 -19.920 ;
        RECT 91.130 -19.970 92.120 -19.920 ;
        RECT 93.010 -19.970 146.400 -19.920 ;
        RECT -45.490 -23.510 146.400 -19.970 ;
        RECT -45.490 -87.220 -43.520 -23.510 ;
      LAYER met1 ;
        RECT -43.520 -87.220 147.150 -23.510 ;
      LAYER met2 ;
        RECT -43.520 -20.700 2.060 50.950 ;
        RECT 2.760 -13.960 7.870 50.950 ;
        RECT 2.760 -14.850 3.050 -13.960 ;
        RECT 3.940 -14.850 6.840 -13.960 ;
        RECT 7.720 -14.850 7.870 -13.960 ;
        RECT 2.760 -18.160 3.140 -14.850 ;
        RECT 3.840 -18.160 6.940 -14.850 ;
        RECT 2.760 -19.050 3.120 -18.160 ;
        RECT 4.010 -18.170 6.940 -18.160 ;
        RECT 7.640 -18.170 7.870 -14.850 ;
        RECT 4.010 -19.050 6.800 -18.170 ;
        RECT 2.760 -19.060 6.800 -19.050 ;
        RECT 7.690 -19.060 7.870 -18.170 ;
        RECT 2.760 -20.680 7.870 -19.060 ;
        RECT 8.570 -13.960 13.580 50.950 ;
        RECT 8.570 -14.850 8.800 -13.960 ;
        RECT 9.690 -14.850 12.590 -13.960 ;
        RECT 13.470 -14.850 13.580 -13.960 ;
        RECT 8.570 -18.160 8.890 -14.850 ;
        RECT 9.590 -18.160 12.690 -14.850 ;
        RECT 8.570 -19.050 8.870 -18.160 ;
        RECT 9.760 -18.170 12.690 -18.160 ;
        RECT 13.390 -18.170 13.580 -14.850 ;
        RECT 9.760 -19.050 12.550 -18.170 ;
        RECT 8.570 -19.060 12.550 -19.050 ;
        RECT 13.440 -19.060 13.580 -18.170 ;
        RECT 8.570 -20.680 13.580 -19.060 ;
        RECT 2.760 -20.700 7.780 -20.680 ;
        RECT -43.520 -21.580 1.970 -20.700 ;
        RECT 2.850 -21.560 7.780 -20.700 ;
        RECT 8.660 -20.690 13.580 -20.680 ;
        RECT 14.280 -13.960 19.360 50.950 ;
        RECT 14.280 -14.850 14.550 -13.960 ;
        RECT 15.440 -14.850 18.340 -13.960 ;
        RECT 19.220 -14.850 19.360 -13.960 ;
        RECT 14.280 -18.160 14.640 -14.850 ;
        RECT 15.340 -18.160 18.440 -14.850 ;
        RECT 14.280 -19.050 14.620 -18.160 ;
        RECT 15.510 -18.170 18.440 -18.160 ;
        RECT 19.140 -18.170 19.360 -14.850 ;
        RECT 15.510 -19.050 18.300 -18.170 ;
        RECT 14.280 -19.060 18.300 -19.050 ;
        RECT 19.190 -19.060 19.360 -18.170 ;
        RECT 14.280 -20.690 19.360 -19.060 ;
        RECT 8.660 -21.560 13.500 -20.690 ;
        RECT 2.850 -21.570 13.500 -21.560 ;
        RECT 14.380 -20.710 19.360 -20.690 ;
        RECT 20.060 -13.960 25.090 50.950 ;
        RECT 20.060 -14.850 20.300 -13.960 ;
        RECT 21.190 -14.850 24.090 -13.960 ;
        RECT 24.970 -14.850 25.090 -13.960 ;
        RECT 20.060 -18.160 20.390 -14.850 ;
        RECT 21.090 -18.160 24.190 -14.850 ;
        RECT 20.060 -19.050 20.370 -18.160 ;
        RECT 21.260 -18.170 24.190 -18.160 ;
        RECT 24.890 -18.170 25.090 -14.850 ;
        RECT 21.260 -19.050 24.050 -18.170 ;
        RECT 20.060 -19.060 24.050 -19.050 ;
        RECT 24.940 -19.060 25.090 -18.170 ;
        RECT 20.060 -20.710 25.090 -19.060 ;
        RECT 25.790 -13.960 30.820 50.950 ;
        RECT 25.790 -14.850 26.050 -13.960 ;
        RECT 26.940 -14.850 29.840 -13.960 ;
        RECT 30.720 -14.850 30.820 -13.960 ;
        RECT 25.790 -18.160 26.140 -14.850 ;
        RECT 26.840 -18.160 29.940 -14.850 ;
        RECT 25.790 -19.050 26.120 -18.160 ;
        RECT 27.010 -18.170 29.940 -18.160 ;
        RECT 30.640 -18.170 30.820 -14.850 ;
        RECT 27.010 -19.050 29.800 -18.170 ;
        RECT 25.790 -19.060 29.800 -19.050 ;
        RECT 30.690 -19.060 30.820 -18.170 ;
        RECT 25.790 -20.710 30.820 -19.060 ;
        RECT 14.380 -21.570 19.280 -20.710 ;
        RECT 2.850 -21.580 19.280 -21.570 ;
        RECT -43.520 -21.590 19.280 -21.580 ;
        RECT 20.160 -21.590 25.030 -20.710 ;
        RECT 25.910 -20.730 30.820 -20.710 ;
        RECT 31.520 -13.960 36.580 50.950 ;
        RECT 31.520 -14.850 31.800 -13.960 ;
        RECT 32.690 -14.850 35.590 -13.960 ;
        RECT 36.470 -14.850 36.580 -13.960 ;
        RECT 31.520 -18.160 31.890 -14.850 ;
        RECT 32.590 -18.160 35.690 -14.850 ;
        RECT 31.520 -19.050 31.870 -18.160 ;
        RECT 32.760 -18.170 35.690 -18.160 ;
        RECT 36.390 -18.170 36.580 -14.850 ;
        RECT 32.760 -19.050 35.550 -18.170 ;
        RECT 31.520 -19.060 35.550 -19.050 ;
        RECT 36.440 -19.060 36.580 -18.170 ;
        RECT 31.520 -20.720 36.580 -19.060 ;
        RECT 37.280 -13.960 42.360 50.950 ;
        RECT 37.280 -14.850 37.550 -13.960 ;
        RECT 38.440 -14.850 41.340 -13.960 ;
        RECT 42.220 -14.850 42.360 -13.960 ;
        RECT 37.280 -18.160 37.640 -14.850 ;
        RECT 38.340 -18.160 41.440 -14.850 ;
        RECT 37.280 -19.050 37.620 -18.160 ;
        RECT 38.510 -18.170 41.440 -18.160 ;
        RECT 42.140 -18.170 42.360 -14.850 ;
        RECT 38.510 -19.050 41.300 -18.170 ;
        RECT 37.280 -19.060 41.300 -19.050 ;
        RECT 42.190 -19.060 42.360 -18.170 ;
        RECT 37.280 -20.710 42.360 -19.060 ;
        RECT 43.060 -13.960 48.090 50.950 ;
        RECT 43.060 -14.850 43.300 -13.960 ;
        RECT 44.190 -14.850 47.090 -13.960 ;
        RECT 47.970 -14.850 48.090 -13.960 ;
        RECT 43.060 -18.160 43.390 -14.850 ;
        RECT 44.090 -18.160 47.190 -14.850 ;
        RECT 43.060 -19.050 43.370 -18.160 ;
        RECT 44.260 -18.170 47.190 -18.160 ;
        RECT 47.890 -18.170 48.090 -14.850 ;
        RECT 44.260 -19.050 47.050 -18.170 ;
        RECT 43.060 -19.060 47.050 -19.050 ;
        RECT 47.940 -19.060 48.090 -18.170 ;
        RECT 43.060 -20.700 48.090 -19.060 ;
        RECT 48.790 -13.960 53.840 50.950 ;
        RECT 48.790 -14.850 49.050 -13.960 ;
        RECT 49.940 -14.850 52.840 -13.960 ;
        RECT 53.720 -14.850 53.840 -13.960 ;
        RECT 48.790 -18.160 49.140 -14.850 ;
        RECT 49.840 -18.160 52.940 -14.850 ;
        RECT 48.790 -19.050 49.120 -18.160 ;
        RECT 50.010 -18.170 52.940 -18.160 ;
        RECT 53.640 -18.170 53.840 -14.850 ;
        RECT 50.010 -19.050 52.800 -18.170 ;
        RECT 48.790 -19.060 52.800 -19.050 ;
        RECT 53.690 -19.060 53.840 -18.170 ;
        RECT 48.790 -20.700 53.840 -19.060 ;
        RECT 43.060 -20.710 48.010 -20.700 ;
        RECT 37.280 -20.720 42.310 -20.710 ;
        RECT 31.520 -20.730 36.510 -20.720 ;
        RECT 25.910 -21.590 30.740 -20.730 ;
        RECT -43.520 -21.610 30.740 -21.590 ;
        RECT 31.620 -21.600 36.510 -20.730 ;
        RECT 37.390 -21.590 42.310 -20.720 ;
        RECT 43.190 -21.580 48.010 -20.710 ;
        RECT 48.890 -20.720 53.840 -20.700 ;
        RECT 54.540 -13.960 59.600 50.950 ;
        RECT 54.540 -14.850 54.800 -13.960 ;
        RECT 55.690 -14.850 58.590 -13.960 ;
        RECT 59.470 -14.850 59.600 -13.960 ;
        RECT 54.540 -18.160 54.890 -14.850 ;
        RECT 55.590 -18.160 58.690 -14.850 ;
        RECT 54.540 -19.050 54.870 -18.160 ;
        RECT 55.760 -18.170 58.690 -18.160 ;
        RECT 59.390 -18.170 59.600 -14.850 ;
        RECT 55.760 -19.050 58.550 -18.170 ;
        RECT 54.540 -19.060 58.550 -19.050 ;
        RECT 59.440 -19.060 59.600 -18.170 ;
        RECT 54.540 -20.700 59.600 -19.060 ;
        RECT 60.300 -13.960 65.330 50.950 ;
        RECT 60.300 -14.850 60.550 -13.960 ;
        RECT 61.440 -14.850 64.340 -13.960 ;
        RECT 65.220 -14.850 65.330 -13.960 ;
        RECT 60.300 -18.160 60.640 -14.850 ;
        RECT 61.340 -18.160 64.440 -14.850 ;
        RECT 60.300 -19.050 60.620 -18.160 ;
        RECT 61.510 -18.170 64.440 -18.160 ;
        RECT 65.140 -18.170 65.330 -14.850 ;
        RECT 61.510 -19.050 64.300 -18.170 ;
        RECT 60.300 -19.060 64.300 -19.050 ;
        RECT 65.190 -19.060 65.330 -18.170 ;
        RECT 60.300 -20.700 65.330 -19.060 ;
        RECT 54.540 -20.720 59.520 -20.700 ;
        RECT 48.890 -21.580 53.780 -20.720 ;
        RECT 43.190 -21.590 53.780 -21.580 ;
        RECT 37.390 -21.600 53.780 -21.590 ;
        RECT 54.660 -21.580 59.520 -20.720 ;
        RECT 60.400 -20.710 65.330 -20.700 ;
        RECT 66.030 -13.960 71.080 50.950 ;
        RECT 66.030 -14.850 66.300 -13.960 ;
        RECT 67.190 -14.850 70.090 -13.960 ;
        RECT 70.970 -14.850 71.080 -13.960 ;
        RECT 66.030 -18.160 66.390 -14.850 ;
        RECT 67.090 -18.160 70.190 -14.850 ;
        RECT 66.030 -19.050 66.370 -18.160 ;
        RECT 67.260 -18.170 70.190 -18.160 ;
        RECT 70.890 -18.170 71.080 -14.850 ;
        RECT 67.260 -19.050 70.050 -18.170 ;
        RECT 66.030 -19.060 70.050 -19.050 ;
        RECT 70.940 -19.060 71.080 -18.170 ;
        RECT 66.030 -20.710 71.080 -19.060 ;
        RECT 60.400 -21.580 65.250 -20.710 ;
        RECT 54.660 -21.590 65.250 -21.580 ;
        RECT 66.130 -20.720 71.080 -20.710 ;
        RECT 71.780 -13.960 76.830 50.950 ;
        RECT 71.780 -14.850 72.050 -13.960 ;
        RECT 72.940 -14.850 75.840 -13.960 ;
        RECT 76.720 -14.850 76.830 -13.960 ;
        RECT 71.780 -18.160 72.140 -14.850 ;
        RECT 72.840 -18.160 75.940 -14.850 ;
        RECT 71.780 -19.050 72.120 -18.160 ;
        RECT 73.010 -18.170 75.940 -18.160 ;
        RECT 76.640 -18.170 76.830 -14.850 ;
        RECT 73.010 -19.050 75.800 -18.170 ;
        RECT 71.780 -19.060 75.800 -19.050 ;
        RECT 76.690 -19.060 76.830 -18.170 ;
        RECT 71.780 -20.720 76.830 -19.060 ;
        RECT 77.530 -13.960 82.600 50.950 ;
        RECT 77.530 -14.850 77.800 -13.960 ;
        RECT 78.690 -14.850 81.590 -13.960 ;
        RECT 82.470 -14.850 82.600 -13.960 ;
        RECT 77.530 -18.160 77.890 -14.850 ;
        RECT 78.590 -18.160 81.690 -14.850 ;
        RECT 77.530 -19.050 77.870 -18.160 ;
        RECT 78.760 -18.170 81.690 -18.160 ;
        RECT 82.390 -18.170 82.600 -14.850 ;
        RECT 78.760 -19.050 81.550 -18.170 ;
        RECT 77.530 -19.060 81.550 -19.050 ;
        RECT 82.440 -19.060 82.600 -18.170 ;
        RECT 77.530 -20.720 82.600 -19.060 ;
        RECT 66.130 -21.590 71.020 -20.720 ;
        RECT 54.660 -21.600 71.020 -21.590 ;
        RECT 71.900 -21.600 76.780 -20.720 ;
        RECT 77.660 -20.740 82.600 -20.720 ;
        RECT 83.300 -13.960 88.350 50.950 ;
        RECT 83.300 -14.850 83.550 -13.960 ;
        RECT 84.440 -14.850 87.340 -13.960 ;
        RECT 88.220 -14.850 88.350 -13.960 ;
        RECT 83.300 -18.160 83.640 -14.850 ;
        RECT 84.340 -18.160 87.440 -14.850 ;
        RECT 83.300 -19.050 83.620 -18.160 ;
        RECT 84.510 -18.170 87.440 -18.160 ;
        RECT 88.140 -18.170 88.350 -14.850 ;
        RECT 84.510 -19.050 87.300 -18.170 ;
        RECT 83.300 -19.060 87.300 -19.050 ;
        RECT 88.190 -19.060 88.350 -18.170 ;
        RECT 83.300 -20.740 88.350 -19.060 ;
        RECT 89.050 -13.960 146.400 50.950 ;
        RECT 89.050 -14.850 89.300 -13.960 ;
        RECT 90.190 -14.850 93.090 -13.960 ;
        RECT 93.970 -14.850 146.400 -13.960 ;
        RECT 89.050 -18.160 89.390 -14.850 ;
        RECT 90.090 -18.160 93.190 -14.850 ;
        RECT 89.050 -19.050 89.370 -18.160 ;
        RECT 90.260 -18.170 93.190 -18.160 ;
        RECT 93.890 -18.170 146.400 -14.850 ;
        RECT 90.260 -19.050 93.050 -18.170 ;
        RECT 89.050 -19.060 93.050 -19.050 ;
        RECT 93.940 -19.060 146.400 -18.170 ;
        RECT 89.050 -20.740 146.400 -19.060 ;
        RECT 77.660 -21.600 82.510 -20.740 ;
        RECT 31.620 -21.610 82.510 -21.600 ;
        RECT -43.520 -21.620 82.510 -21.610 ;
        RECT 83.390 -21.620 88.260 -20.740 ;
        RECT 89.140 -21.620 146.400 -20.740 ;
        RECT -43.520 -23.510 146.400 -21.620 ;
      LAYER met2 ;
        RECT -43.520 -87.220 147.150 -23.510 ;
      LAYER met3 ;
        RECT 100.780 49.940 146.400 50.950 ;
        RECT -42.410 49.930 62.290 49.940 ;
        RECT 63.490 49.930 146.400 49.940 ;
        RECT -42.410 49.880 146.400 49.930 ;
        RECT -43.520 -5.640 146.400 49.880 ;
        RECT -43.520 -6.800 5.530 -5.640 ;
        RECT 6.690 -5.670 146.400 -5.640 ;
        RECT 100.880 -6.770 146.400 -5.670 ;
        RECT 6.690 -6.800 146.400 -6.770 ;
        RECT -43.520 -6.910 146.400 -6.800 ;
        RECT -43.520 -8.070 11.280 -6.910 ;
        RECT 12.440 -6.940 146.400 -6.910 ;
        RECT 100.880 -8.040 146.400 -6.940 ;
        RECT 12.440 -8.070 146.400 -8.040 ;
        RECT -43.520 -8.280 146.400 -8.070 ;
        RECT -43.520 -9.440 17.080 -8.280 ;
        RECT 18.240 -8.310 146.400 -8.280 ;
        RECT 100.880 -9.410 146.400 -8.310 ;
        RECT 18.240 -9.440 146.400 -9.410 ;
        RECT -43.520 -9.450 146.400 -9.440 ;
        RECT -43.520 -10.610 22.780 -9.450 ;
        RECT 23.940 -9.480 146.400 -9.450 ;
        RECT 100.880 -10.580 146.400 -9.480 ;
        RECT 23.940 -10.610 146.400 -10.580 ;
        RECT -43.520 -10.700 146.400 -10.610 ;
        RECT -43.520 -11.860 28.530 -10.700 ;
        RECT 29.690 -10.730 146.400 -10.700 ;
        RECT 100.880 -11.830 146.400 -10.730 ;
        RECT 29.690 -11.860 146.400 -11.830 ;
        RECT -43.520 -12.150 146.400 -11.860 ;
        RECT -43.520 -13.310 34.280 -12.150 ;
        RECT 35.440 -12.180 146.400 -12.150 ;
        RECT 100.880 -13.280 146.400 -12.180 ;
        RECT 35.440 -13.310 146.400 -13.280 ;
        RECT -43.520 -13.350 146.400 -13.310 ;
        RECT -43.520 -14.550 40.000 -13.350 ;
        RECT 41.200 -13.400 146.400 -13.350 ;
        RECT 41.200 -14.550 45.780 -14.500 ;
        RECT -43.520 -15.410 45.780 -14.550 ;
        RECT 46.940 -15.410 51.530 -15.380 ;
        RECT -43.520 -16.240 51.530 -15.410 ;
        RECT 52.690 -16.240 57.280 -16.210 ;
        RECT -43.520 -17.020 57.280 -16.240 ;
        RECT 58.440 -17.020 63.030 -16.990 ;
        RECT -43.520 -17.880 63.030 -17.020 ;
        RECT 64.190 -17.880 68.780 -17.850 ;
        RECT -43.520 -18.680 68.780 -17.880 ;
        RECT 69.940 -18.680 74.530 -18.650 ;
        RECT -43.520 -19.480 74.530 -18.680 ;
        RECT 75.690 -19.480 80.280 -19.450 ;
        RECT -43.520 -19.850 80.280 -19.480 ;
        RECT -43.520 -19.900 -0.800 -19.850 ;
        RECT 0.400 -20.130 80.280 -19.850 ;
        RECT 100.880 -20.100 146.400 -13.400 ;
        RECT 81.440 -20.110 146.400 -20.100 ;
        RECT 81.440 -20.130 86.030 -20.110 ;
        RECT -43.520 -21.070 -42.230 -21.000 ;
        RECT -41.070 -21.050 -0.800 -21.000 ;
        RECT 0.400 -21.050 86.030 -20.130 ;
        RECT 87.190 -20.140 146.400 -20.110 ;
        RECT -41.070 -21.070 -0.750 -21.050 ;
        RECT -43.520 -23.510 -0.750 -21.070 ;
        RECT 0.350 -21.270 86.030 -21.050 ;
        RECT 87.190 -21.270 91.780 -21.240 ;
        RECT 0.350 -22.160 91.780 -21.270 ;
        RECT 100.880 -22.130 146.400 -20.140 ;
        RECT 92.940 -22.160 146.400 -22.130 ;
        RECT 0.350 -22.740 146.400 -22.160 ;
        RECT 0.350 -22.750 88.250 -22.740 ;
        RECT 0.350 -22.800 7.660 -22.750 ;
        RECT 8.860 -22.760 88.250 -22.750 ;
        RECT 0.350 -22.810 7.650 -22.800 ;
        RECT 8.860 -22.810 19.150 -22.760 ;
        RECT 20.350 -22.770 53.550 -22.760 ;
        RECT 20.350 -22.810 30.580 -22.770 ;
        RECT 31.780 -22.780 53.550 -22.770 ;
        RECT 31.780 -22.810 42.150 -22.780 ;
        RECT 43.350 -22.810 53.550 -22.780 ;
        RECT 54.750 -22.810 65.230 -22.760 ;
        RECT 66.430 -22.810 76.680 -22.760 ;
        RECT 77.880 -22.790 88.250 -22.760 ;
        RECT 77.880 -22.810 88.240 -22.790 ;
        RECT 89.450 -23.510 146.400 -22.740 ;
      LAYER met3 ;
        RECT -43.520 -87.220 147.150 -23.510 ;
  END
END Integrated_bitcell_with_dummy_cells
END LIBRARY

